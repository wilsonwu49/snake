library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity currscore_rom is
  port (
    x     : in  std_logic_vector(4 downto 0);
    y     : in  std_logic_vector(3 downto 0);
    pixel : out std_logic_vector(5 downto 0)
  );
end entity;


architecture synth of currscore_rom is
  signal addr : unsigned(8 downto 0);
  
  attribute syn_ramstyle : string;
	attribute syn_ramstyle of pixel : signal is "registers" ;
begin
  addr <= resize((unsigned(y) * 32) + unsigned(x), 9);
  process(addr)
  begin
    case addr is
      when 0 => pixel <= "111111";
      when 1 => pixel <= "111111";
      when 2 => pixel <= "111111";
      when 3 => pixel <= "111111";
      when 4 => pixel <= "111111";
      when 5 => pixel <= "111111";
      when 6 => pixel <= "111111";
      when 7 => pixel <= "111111";
      when 8 => pixel <= "111111";
      when 9 => pixel <= "111111";
      when 10 => pixel <= "111111";
      when 11 => pixel <= "111111";
      when 12 => pixel <= "111111";
      when 13 => pixel <= "111111";
      when 14 => pixel <= "111111";
      when 15 => pixel <= "111111";
      when 16 => pixel <= "111111";
      when 17 => pixel <= "111111";
      when 18 => pixel <= "111111";
      when 19 => pixel <= "111111";
      when 20 => pixel <= "111111";
      when 21 => pixel <= "111111";
      when 22 => pixel <= "111111";
      when 23 => pixel <= "111111";
      when 24 => pixel <= "111111";
      when 25 => pixel <= "111111";
      when 26 => pixel <= "111111";
      when 27 => pixel <= "111111";
      when 28 => pixel <= "111111";
      when 29 => pixel <= "111111";
      when 30 => pixel <= "111111";
      when 31 => pixel <= "111111";
      when 32 => pixel <= "111111";
      when 33 => pixel <= "111111";
      when 34 => pixel <= "111111";
      when 35 => pixel <= "111111";
      when 36 => pixel <= "111111";
      when 37 => pixel <= "111111";
      when 38 => pixel <= "111111";
      when 39 => pixel <= "111111";
      when 40 => pixel <= "111111";
      when 41 => pixel <= "111111";
      when 42 => pixel <= "111111";
      when 43 => pixel <= "111111";
      when 44 => pixel <= "111111";
      when 45 => pixel <= "111111";
      when 46 => pixel <= "111111";
      when 47 => pixel <= "111111";
      when 48 => pixel <= "111111";
      when 49 => pixel <= "111111";
      when 50 => pixel <= "111111";
      when 51 => pixel <= "111111";
      when 52 => pixel <= "111111";
      when 53 => pixel <= "111111";
      when 54 => pixel <= "111111";
      when 55 => pixel <= "111111";
      when 56 => pixel <= "111111";
      when 57 => pixel <= "111111";
      when 58 => pixel <= "111111";
      when 59 => pixel <= "111111";
      when 60 => pixel <= "111111";
      when 61 => pixel <= "111111";
      when 62 => pixel <= "111111";
      when 63 => pixel <= "111111";
      when 64 => pixel <= "111111";
      when 65 => pixel <= "111111";
      when 66 => pixel <= "111111";
      when 67 => pixel <= "111111";
      when 68 => pixel <= "111111";
      when 69 => pixel <= "111111";
      when 70 => pixel <= "000000";
      when 71 => pixel <= "000000";
      when 72 => pixel <= "111111";
      when 73 => pixel <= "111111";
      when 74 => pixel <= "000000";
      when 75 => pixel <= "111111";
      when 76 => pixel <= "111111";
      when 77 => pixel <= "000000";
      when 78 => pixel <= "111111";
      when 79 => pixel <= "000000";
      when 80 => pixel <= "000000";
      when 81 => pixel <= "000000";
      when 82 => pixel <= "111111";
      when 83 => pixel <= "111111";
      when 84 => pixel <= "000000";
      when 85 => pixel <= "000000";
      when 86 => pixel <= "000000";
      when 87 => pixel <= "111111";
      when 88 => pixel <= "111111";
      when 89 => pixel <= "111111";
      when 90 => pixel <= "111111";
      when 91 => pixel <= "111111";
      when 92 => pixel <= "111111";
      when 93 => pixel <= "111111";
      when 94 => pixel <= "111111";
      when 95 => pixel <= "111111";
      when 96 => pixel <= "111111";
      when 97 => pixel <= "111111";
      when 98 => pixel <= "111111";
      when 99 => pixel <= "111111";
      when 100 => pixel <= "111111";
      when 101 => pixel <= "000000";
      when 102 => pixel <= "111111";
      when 103 => pixel <= "111111";
      when 104 => pixel <= "000000";
      when 105 => pixel <= "111111";
      when 106 => pixel <= "000000";
      when 107 => pixel <= "111111";
      when 108 => pixel <= "111111";
      when 109 => pixel <= "000000";
      when 110 => pixel <= "111111";
      when 111 => pixel <= "000000";
      when 112 => pixel <= "111111";
      when 113 => pixel <= "111111";
      when 114 => pixel <= "000000";
      when 115 => pixel <= "111111";
      when 116 => pixel <= "000000";
      when 117 => pixel <= "111111";
      when 118 => pixel <= "111111";
      when 119 => pixel <= "000000";
      when 120 => pixel <= "111111";
      when 121 => pixel <= "111111";
      when 122 => pixel <= "111111";
      when 123 => pixel <= "111111";
      when 124 => pixel <= "111111";
      when 125 => pixel <= "111111";
      when 126 => pixel <= "111111";
      when 127 => pixel <= "111111";
      when 128 => pixel <= "111111";
      when 129 => pixel <= "111111";
      when 130 => pixel <= "111111";
      when 131 => pixel <= "111111";
      when 132 => pixel <= "111111";
      when 133 => pixel <= "000000";
      when 134 => pixel <= "111111";
      when 135 => pixel <= "111111";
      when 136 => pixel <= "111111";
      when 137 => pixel <= "111111";
      when 138 => pixel <= "000000";
      when 139 => pixel <= "111111";
      when 140 => pixel <= "111111";
      when 141 => pixel <= "000000";
      when 142 => pixel <= "111111";
      when 143 => pixel <= "000000";
      when 144 => pixel <= "000000";
      when 145 => pixel <= "000000";
      when 146 => pixel <= "111111";
      when 147 => pixel <= "111111";
      when 148 => pixel <= "000000";
      when 149 => pixel <= "000000";
      when 150 => pixel <= "000000";
      when 151 => pixel <= "111111";
      when 152 => pixel <= "111111";
      when 153 => pixel <= "111111";
      when 154 => pixel <= "111111";
      when 155 => pixel <= "111111";
      when 156 => pixel <= "111111";
      when 157 => pixel <= "111111";
      when 158 => pixel <= "111111";
      when 159 => pixel <= "111111";
      when 160 => pixel <= "111111";
      when 161 => pixel <= "111111";
      when 162 => pixel <= "111111";
      when 163 => pixel <= "111111";
      when 164 => pixel <= "111111";
      when 165 => pixel <= "000000";
      when 166 => pixel <= "111111";
      when 167 => pixel <= "111111";
      when 168 => pixel <= "000000";
      when 169 => pixel <= "111111";
      when 170 => pixel <= "000000";
      when 171 => pixel <= "111111";
      when 172 => pixel <= "111111";
      when 173 => pixel <= "000000";
      when 174 => pixel <= "111111";
      when 175 => pixel <= "000000";
      when 176 => pixel <= "111111";
      when 177 => pixel <= "000000";
      when 178 => pixel <= "111111";
      when 179 => pixel <= "111111";
      when 180 => pixel <= "000000";
      when 181 => pixel <= "111111";
      when 182 => pixel <= "000000";
      when 183 => pixel <= "111111";
      when 184 => pixel <= "111111";
      when 185 => pixel <= "111111";
      when 186 => pixel <= "111111";
      when 187 => pixel <= "111111";
      when 188 => pixel <= "111111";
      when 189 => pixel <= "111111";
      when 190 => pixel <= "111111";
      when 191 => pixel <= "111111";
      when 192 => pixel <= "111111";
      when 193 => pixel <= "111111";
      when 194 => pixel <= "111111";
      when 195 => pixel <= "111111";
      when 196 => pixel <= "111111";
      when 197 => pixel <= "111111";
      when 198 => pixel <= "000000";
      when 199 => pixel <= "000000";
      when 200 => pixel <= "111111";
      when 201 => pixel <= "111111";
      when 202 => pixel <= "111111";
      when 203 => pixel <= "000000";
      when 204 => pixel <= "000000";
      when 205 => pixel <= "111111";
      when 206 => pixel <= "111111";
      when 207 => pixel <= "000000";
      when 208 => pixel <= "111111";
      when 209 => pixel <= "111111";
      when 210 => pixel <= "000000";
      when 211 => pixel <= "111111";
      when 212 => pixel <= "000000";
      when 213 => pixel <= "111111";
      when 214 => pixel <= "111111";
      when 215 => pixel <= "000000";
      when 216 => pixel <= "111111";
      when 217 => pixel <= "111111";
      when 218 => pixel <= "000000";
      when 219 => pixel <= "111111";
      when 220 => pixel <= "111111";
      when 221 => pixel <= "111111";
      when 222 => pixel <= "111111";
      when 223 => pixel <= "111111";
      when 224 => pixel <= "111111";
      when 225 => pixel <= "111111";
      when 226 => pixel <= "111111";
      when 227 => pixel <= "111111";
      when 228 => pixel <= "111111";
      when 229 => pixel <= "111111";
      when 230 => pixel <= "111111";
      when 231 => pixel <= "111111";
      when 232 => pixel <= "111111";
      when 233 => pixel <= "111111";
      when 234 => pixel <= "111111";
      when 235 => pixel <= "111111";
      when 236 => pixel <= "111111";
      when 237 => pixel <= "111111";
      when 238 => pixel <= "111111";
      when 239 => pixel <= "111111";
      when 240 => pixel <= "111111";
      when 241 => pixel <= "111111";
      when 242 => pixel <= "111111";
      when 243 => pixel <= "111111";
      when 244 => pixel <= "111111";
      when 245 => pixel <= "111111";
      when 246 => pixel <= "111111";
      when 247 => pixel <= "111111";
      when 248 => pixel <= "111111";
      when 249 => pixel <= "111111";
      when 250 => pixel <= "111111";
      when 251 => pixel <= "111111";
      when 252 => pixel <= "111111";
      when 253 => pixel <= "111111";
      when 254 => pixel <= "111111";
      when 255 => pixel <= "111111";
      when 256 => pixel <= "111111";
      when 257 => pixel <= "111111";
      when 258 => pixel <= "111111";
      when 259 => pixel <= "111111";
      when 260 => pixel <= "111111";
      when 261 => pixel <= "111111";
      when 262 => pixel <= "111111";
      when 263 => pixel <= "111111";
      when 264 => pixel <= "111111";
      when 265 => pixel <= "111111";
      when 266 => pixel <= "111111";
      when 267 => pixel <= "111111";
      when 268 => pixel <= "111111";
      when 269 => pixel <= "111111";
      when 270 => pixel <= "111111";
      when 271 => pixel <= "111111";
      when 272 => pixel <= "111111";
      when 273 => pixel <= "111111";
      when 274 => pixel <= "111111";
      when 275 => pixel <= "111111";
      when 276 => pixel <= "111111";
      when 277 => pixel <= "111111";
      when 278 => pixel <= "111111";
      when 279 => pixel <= "111111";
      when 280 => pixel <= "111111";
      when 281 => pixel <= "111111";
      when 282 => pixel <= "111111";
      when 283 => pixel <= "111111";
      when 284 => pixel <= "111111";
      when 285 => pixel <= "111111";
      when 286 => pixel <= "111111";
      when 287 => pixel <= "111111";
      when 288 => pixel <= "111111";
      when 289 => pixel <= "111111";
      when 290 => pixel <= "111111";
      when 291 => pixel <= "111111";
      when 292 => pixel <= "111111";
      when 293 => pixel <= "000000";
      when 294 => pixel <= "000000";
      when 295 => pixel <= "000000";
      when 296 => pixel <= "111111";
      when 297 => pixel <= "111111";
      when 298 => pixel <= "000000";
      when 299 => pixel <= "000000";
      when 300 => pixel <= "111111";
      when 301 => pixel <= "111111";
      when 302 => pixel <= "111111";
      when 303 => pixel <= "000000";
      when 304 => pixel <= "000000";
      when 305 => pixel <= "111111";
      when 306 => pixel <= "111111";
      when 307 => pixel <= "000000";
      when 308 => pixel <= "000000";
      when 309 => pixel <= "000000";
      when 310 => pixel <= "111111";
      when 311 => pixel <= "111111";
      when 312 => pixel <= "000000";
      when 313 => pixel <= "000000";
      when 314 => pixel <= "000000";
      when 315 => pixel <= "000000";
      when 316 => pixel <= "111111";
      when 317 => pixel <= "111111";
      when 318 => pixel <= "111111";
      when 319 => pixel <= "111111";
      when 320 => pixel <= "111111";
      when 321 => pixel <= "111111";
      when 322 => pixel <= "111111";
      when 323 => pixel <= "111111";
      when 324 => pixel <= "000000";
      when 325 => pixel <= "111111";
      when 326 => pixel <= "111111";
      when 327 => pixel <= "111111";
      when 328 => pixel <= "111111";
      when 329 => pixel <= "000000";
      when 330 => pixel <= "111111";
      when 331 => pixel <= "111111";
      when 332 => pixel <= "000000";
      when 333 => pixel <= "111111";
      when 334 => pixel <= "000000";
      when 335 => pixel <= "111111";
      when 336 => pixel <= "111111";
      when 337 => pixel <= "000000";
      when 338 => pixel <= "111111";
      when 339 => pixel <= "000000";
      when 340 => pixel <= "111111";
      when 341 => pixel <= "111111";
      when 342 => pixel <= "000000";
      when 343 => pixel <= "111111";
      when 344 => pixel <= "000000";
      when 345 => pixel <= "111111";
      when 346 => pixel <= "111111";
      when 347 => pixel <= "111111";
      when 348 => pixel <= "111111";
      when 349 => pixel <= "111111";
      when 350 => pixel <= "111111";
      when 351 => pixel <= "111111";
      when 352 => pixel <= "111111";
      when 353 => pixel <= "111111";
      when 354 => pixel <= "111111";
      when 355 => pixel <= "111111";
      when 356 => pixel <= "111111";
      when 357 => pixel <= "000000";
      when 358 => pixel <= "000000";
      when 359 => pixel <= "111111";
      when 360 => pixel <= "111111";
      when 361 => pixel <= "000000";
      when 362 => pixel <= "111111";
      when 363 => pixel <= "111111";
      when 364 => pixel <= "111111";
      when 365 => pixel <= "111111";
      when 366 => pixel <= "000000";
      when 367 => pixel <= "111111";
      when 368 => pixel <= "111111";
      when 369 => pixel <= "000000";
      when 370 => pixel <= "111111";
      when 371 => pixel <= "000000";
      when 372 => pixel <= "000000";
      when 373 => pixel <= "000000";
      when 374 => pixel <= "111111";
      when 375 => pixel <= "111111";
      when 376 => pixel <= "000000";
      when 377 => pixel <= "000000";
      when 378 => pixel <= "000000";
      when 379 => pixel <= "111111";
      when 380 => pixel <= "111111";
      when 381 => pixel <= "111111";
      when 382 => pixel <= "111111";
      when 383 => pixel <= "111111";
      when 384 => pixel <= "111111";
      when 385 => pixel <= "111111";
      when 386 => pixel <= "111111";
      when 387 => pixel <= "111111";
      when 388 => pixel <= "111111";
      when 389 => pixel <= "111111";
      when 390 => pixel <= "111111";
      when 391 => pixel <= "000000";
      when 392 => pixel <= "111111";
      when 393 => pixel <= "000000";
      when 394 => pixel <= "111111";
      when 395 => pixel <= "111111";
      when 396 => pixel <= "000000";
      when 397 => pixel <= "111111";
      when 398 => pixel <= "000000";
      when 399 => pixel <= "111111";
      when 400 => pixel <= "111111";
      when 401 => pixel <= "000000";
      when 402 => pixel <= "111111";
      when 403 => pixel <= "000000";
      when 404 => pixel <= "111111";
      when 405 => pixel <= "000000";
      when 406 => pixel <= "111111";
      when 407 => pixel <= "111111";
      when 408 => pixel <= "000000";
      when 409 => pixel <= "111111";
      when 410 => pixel <= "111111";
      when 411 => pixel <= "111111";
      when 412 => pixel <= "111111";
      when 413 => pixel <= "111111";
      when 414 => pixel <= "111111";
      when 415 => pixel <= "111111";
      when 416 => pixel <= "111111";
      when 417 => pixel <= "111111";
      when 418 => pixel <= "111111";
      when 419 => pixel <= "111111";
      when 420 => pixel <= "000000";
      when 421 => pixel <= "000000";
      when 422 => pixel <= "000000";
      when 423 => pixel <= "111111";
      when 424 => pixel <= "111111";
      when 425 => pixel <= "111111";
      when 426 => pixel <= "000000";
      when 427 => pixel <= "000000";
      when 428 => pixel <= "111111";
      when 429 => pixel <= "111111";
      when 430 => pixel <= "111111";
      when 431 => pixel <= "000000";
      when 432 => pixel <= "000000";
      when 433 => pixel <= "111111";
      when 434 => pixel <= "111111";
      when 435 => pixel <= "000000";
      when 436 => pixel <= "111111";
      when 437 => pixel <= "111111";
      when 438 => pixel <= "000000";
      when 439 => pixel <= "111111";
      when 440 => pixel <= "000000";
      when 441 => pixel <= "000000";
      when 442 => pixel <= "000000";
      when 443 => pixel <= "000000";
      when 444 => pixel <= "111111";
      when 445 => pixel <= "111111";
      when 446 => pixel <= "111111";
      when 447 => pixel <= "111111";
      when 448 => pixel <= "111111";
      when 449 => pixel <= "111111";
      when 450 => pixel <= "111111";
      when 451 => pixel <= "111111";
      when 452 => pixel <= "111111";
      when 453 => pixel <= "111111";
      when 454 => pixel <= "111111";
      when 455 => pixel <= "111111";
      when 456 => pixel <= "111111";
      when 457 => pixel <= "111111";
      when 458 => pixel <= "111111";
      when 459 => pixel <= "111111";
      when 460 => pixel <= "111111";
      when 461 => pixel <= "111111";
      when 462 => pixel <= "111111";
      when 463 => pixel <= "111111";
      when 464 => pixel <= "111111";
      when 465 => pixel <= "111111";
      when 466 => pixel <= "111111";
      when 467 => pixel <= "111111";
      when 468 => pixel <= "111111";
      when 469 => pixel <= "111111";
      when 470 => pixel <= "111111";
      when 471 => pixel <= "111111";
      when 472 => pixel <= "111111";
      when 473 => pixel <= "111111";
      when 474 => pixel <= "111111";
      when 475 => pixel <= "111111";
      when 476 => pixel <= "111111";
      when 477 => pixel <= "111111";
      when 478 => pixel <= "111111";
      when 479 => pixel <= "111111";
      when 480 => pixel <= "111111";
      when 481 => pixel <= "111111";
      when 482 => pixel <= "111111";
      when 483 => pixel <= "111111";
      when 484 => pixel <= "111111";
      when 485 => pixel <= "111111";
      when 486 => pixel <= "111111";
      when 487 => pixel <= "111111";
      when 488 => pixel <= "111111";
      when 489 => pixel <= "111111";
      when 490 => pixel <= "111111";
      when 491 => pixel <= "111111";
      when 492 => pixel <= "111111";
      when 493 => pixel <= "111111";
      when 494 => pixel <= "111111";
      when 495 => pixel <= "111111";
      when 496 => pixel <= "111111";
      when 497 => pixel <= "111111";
      when 498 => pixel <= "111111";
      when 499 => pixel <= "111111";
      when 500 => pixel <= "111111";
      when 501 => pixel <= "111111";
      when 502 => pixel <= "111111";
      when 503 => pixel <= "111111";
      when 504 => pixel <= "111111";
      when 505 => pixel <= "111111";
      when 506 => pixel <= "111111";
      when 507 => pixel <= "111111";
      when 508 => pixel <= "111111";
      when 509 => pixel <= "111111";
      when 510 => pixel <= "111111";
      when 511 => pixel <= "111111";
      when others => pixel <= (others => '0');
    end case;
  end process;
end;

