library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity gameover_rom is
  port (
    x     : in  std_logic_vector(7 downto 0);
    y     : in  std_logic_vector(6 downto 0);
    pixel : out std_logic_vector(5 downto 0)
  );
end entity;

architecture synth of gameover_rom is
  signal addr : unsigned(14 downto 0);
begin
  addr <= (unsigned(y) * 8d"160") + unsigned(x);
  process(addr)
  begin
    case addr is
      when 0 => pixel <= "000000";
      when 1 => pixel <= "000000";
      when 2 => pixel <= "000000";
      when 3 => pixel <= "000000";
      when 4 => pixel <= "000000";
      when 5 => pixel <= "000000";
      when 6 => pixel <= "000000";
      when 7 => pixel <= "000000";
      when 8 => pixel <= "000000";
      when 9 => pixel <= "000000";
      when 10 => pixel <= "000000";
      when 11 => pixel <= "000000";
      when 12 => pixel <= "000000";
      when 13 => pixel <= "000000";
      when 14 => pixel <= "000000";
      when 15 => pixel <= "000000";
      when 16 => pixel <= "000000";
      when 17 => pixel <= "000000";
      when 18 => pixel <= "000000";
      when 19 => pixel <= "000000";
      when 20 => pixel <= "000000";
      when 21 => pixel <= "000000";
      when 22 => pixel <= "000000";
      when 23 => pixel <= "000000";
      when 24 => pixel <= "000000";
      when 25 => pixel <= "000000";
      when 26 => pixel <= "000000";
      when 27 => pixel <= "000000";
      when 28 => pixel <= "000000";
      when 29 => pixel <= "000000";
      when 30 => pixel <= "000000";
      when 31 => pixel <= "000000";
      when 32 => pixel <= "000000";
      when 33 => pixel <= "000000";
      when 34 => pixel <= "000000";
      when 35 => pixel <= "000000";
      when 36 => pixel <= "000000";
      when 37 => pixel <= "000000";
      when 38 => pixel <= "000000";
      when 39 => pixel <= "000000";
      when 40 => pixel <= "000000";
      when 41 => pixel <= "000000";
      when 42 => pixel <= "000000";
      when 43 => pixel <= "000000";
      when 44 => pixel <= "000000";
      when 45 => pixel <= "000000";
      when 46 => pixel <= "000000";
      when 47 => pixel <= "000000";
      when 48 => pixel <= "000000";
      when 49 => pixel <= "000000";
      when 50 => pixel <= "000000";
      when 51 => pixel <= "000000";
      when 52 => pixel <= "000000";
      when 53 => pixel <= "000000";
      when 54 => pixel <= "000000";
      when 55 => pixel <= "000000";
      when 56 => pixel <= "000000";
      when 57 => pixel <= "000000";
      when 58 => pixel <= "000000";
      when 59 => pixel <= "000000";
      when 60 => pixel <= "000000";
      when 61 => pixel <= "000000";
      when 62 => pixel <= "000000";
      when 63 => pixel <= "000000";
      when 64 => pixel <= "000000";
      when 65 => pixel <= "000000";
      when 66 => pixel <= "000000";
      when 67 => pixel <= "000000";
      when 68 => pixel <= "000000";
      when 69 => pixel <= "000000";
      when 70 => pixel <= "000000";
      when 71 => pixel <= "000000";
      when 72 => pixel <= "000000";
      when 73 => pixel <= "000000";
      when 74 => pixel <= "000000";
      when 75 => pixel <= "000000";
      when 76 => pixel <= "000000";
      when 77 => pixel <= "000000";
      when 78 => pixel <= "000000";
      when 79 => pixel <= "000000";
      when 80 => pixel <= "000000";
      when 81 => pixel <= "000000";
      when 82 => pixel <= "000000";
      when 83 => pixel <= "000000";
      when 84 => pixel <= "000000";
      when 85 => pixel <= "000000";
      when 86 => pixel <= "000000";
      when 87 => pixel <= "000000";
      when 88 => pixel <= "000000";
      when 89 => pixel <= "000000";
      when 90 => pixel <= "000000";
      when 91 => pixel <= "000000";
      when 92 => pixel <= "000000";
      when 93 => pixel <= "000000";
      when 94 => pixel <= "000000";
      when 95 => pixel <= "000000";
      when 96 => pixel <= "000000";
      when 97 => pixel <= "000000";
      when 98 => pixel <= "000000";
      when 99 => pixel <= "000000";
      when 100 => pixel <= "000000";
      when 101 => pixel <= "000000";
      when 102 => pixel <= "000000";
      when 103 => pixel <= "000000";
      when 104 => pixel <= "000000";
      when 105 => pixel <= "000000";
      when 106 => pixel <= "000000";
      when 107 => pixel <= "000000";
      when 108 => pixel <= "000000";
      when 109 => pixel <= "000000";
      when 110 => pixel <= "000000";
      when 111 => pixel <= "000000";
      when 112 => pixel <= "000000";
      when 113 => pixel <= "000000";
      when 114 => pixel <= "000000";
      when 115 => pixel <= "000000";
      when 116 => pixel <= "000000";
      when 117 => pixel <= "000000";
      when 118 => pixel <= "000000";
      when 119 => pixel <= "000000";
      when 120 => pixel <= "000000";
      when 121 => pixel <= "000000";
      when 122 => pixel <= "000000";
      when 123 => pixel <= "000000";
      when 124 => pixel <= "000000";
      when 125 => pixel <= "000000";
      when 126 => pixel <= "000000";
      when 127 => pixel <= "000000";
      when 128 => pixel <= "000000";
      when 129 => pixel <= "000000";
      when 130 => pixel <= "000000";
      when 131 => pixel <= "000000";
      when 132 => pixel <= "000000";
      when 133 => pixel <= "000000";
      when 134 => pixel <= "000000";
      when 135 => pixel <= "000000";
      when 136 => pixel <= "000000";
      when 137 => pixel <= "000000";
      when 138 => pixel <= "000000";
      when 139 => pixel <= "000000";
      when 140 => pixel <= "000000";
      when 141 => pixel <= "000000";
      when 142 => pixel <= "000000";
      when 143 => pixel <= "000000";
      when 144 => pixel <= "000000";
      when 145 => pixel <= "000000";
      when 146 => pixel <= "000000";
      when 147 => pixel <= "000000";
      when 148 => pixel <= "000000";
      when 149 => pixel <= "000000";
      when 150 => pixel <= "000000";
      when 151 => pixel <= "000000";
      when 152 => pixel <= "000000";
      when 153 => pixel <= "000000";
      when 154 => pixel <= "000000";
      when 155 => pixel <= "000000";
      when 156 => pixel <= "000000";
      when 157 => pixel <= "000000";
      when 158 => pixel <= "000000";
      when 159 => pixel <= "000000";
      when 160 => pixel <= "000000";
      when 161 => pixel <= "000000";
      when 162 => pixel <= "000000";
      when 163 => pixel <= "000000";
      when 164 => pixel <= "000000";
      when 165 => pixel <= "000000";
      when 166 => pixel <= "000000";
      when 167 => pixel <= "000000";
      when 168 => pixel <= "000000";
      when 169 => pixel <= "000000";
      when 170 => pixel <= "000000";
      when 171 => pixel <= "000000";
      when 172 => pixel <= "000000";
      when 173 => pixel <= "000000";
      when 174 => pixel <= "000000";
      when 175 => pixel <= "000000";
      when 176 => pixel <= "000000";
      when 177 => pixel <= "000000";
      when 178 => pixel <= "000000";
      when 179 => pixel <= "000000";
      when 180 => pixel <= "000000";
      when 181 => pixel <= "000000";
      when 182 => pixel <= "000000";
      when 183 => pixel <= "000000";
      when 184 => pixel <= "000000";
      when 185 => pixel <= "000000";
      when 186 => pixel <= "000000";
      when 187 => pixel <= "000000";
      when 188 => pixel <= "000000";
      when 189 => pixel <= "000000";
      when 190 => pixel <= "000000";
      when 191 => pixel <= "000000";
      when 192 => pixel <= "000000";
      when 193 => pixel <= "000000";
      when 194 => pixel <= "000000";
      when 195 => pixel <= "000000";
      when 196 => pixel <= "000000";
      when 197 => pixel <= "000000";
      when 198 => pixel <= "000000";
      when 199 => pixel <= "000000";
      when 200 => pixel <= "000000";
      when 201 => pixel <= "000000";
      when 202 => pixel <= "000000";
      when 203 => pixel <= "000000";
      when 204 => pixel <= "000000";
      when 205 => pixel <= "000000";
      when 206 => pixel <= "000000";
      when 207 => pixel <= "000000";
      when 208 => pixel <= "000000";
      when 209 => pixel <= "000000";
      when 210 => pixel <= "000000";
      when 211 => pixel <= "000000";
      when 212 => pixel <= "000000";
      when 213 => pixel <= "000000";
      when 214 => pixel <= "000000";
      when 215 => pixel <= "000000";
      when 216 => pixel <= "000000";
      when 217 => pixel <= "000000";
      when 218 => pixel <= "000000";
      when 219 => pixel <= "000000";
      when 220 => pixel <= "000000";
      when 221 => pixel <= "000000";
      when 222 => pixel <= "000000";
      when 223 => pixel <= "000000";
      when 224 => pixel <= "000000";
      when 225 => pixel <= "000000";
      when 226 => pixel <= "000000";
      when 227 => pixel <= "000000";
      when 228 => pixel <= "000000";
      when 229 => pixel <= "000000";
      when 230 => pixel <= "000000";
      when 231 => pixel <= "000000";
      when 232 => pixel <= "000000";
      when 233 => pixel <= "000000";
      when 234 => pixel <= "000000";
      when 235 => pixel <= "000000";
      when 236 => pixel <= "000000";
      when 237 => pixel <= "000000";
      when 238 => pixel <= "000000";
      when 239 => pixel <= "000000";
      when 240 => pixel <= "000000";
      when 241 => pixel <= "000000";
      when 242 => pixel <= "000000";
      when 243 => pixel <= "000000";
      when 244 => pixel <= "000000";
      when 245 => pixel <= "000000";
      when 246 => pixel <= "000000";
      when 247 => pixel <= "000000";
      when 248 => pixel <= "000000";
      when 249 => pixel <= "000000";
      when 250 => pixel <= "000000";
      when 251 => pixel <= "000000";
      when 252 => pixel <= "000000";
      when 253 => pixel <= "000000";
      when 254 => pixel <= "000000";
      when 255 => pixel <= "000000";
      when 256 => pixel <= "000000";
      when 257 => pixel <= "000000";
      when 258 => pixel <= "000000";
      when 259 => pixel <= "000000";
      when 260 => pixel <= "000000";
      when 261 => pixel <= "000000";
      when 262 => pixel <= "000000";
      when 263 => pixel <= "000000";
      when 264 => pixel <= "000000";
      when 265 => pixel <= "000000";
      when 266 => pixel <= "000000";
      when 267 => pixel <= "000000";
      when 268 => pixel <= "000000";
      when 269 => pixel <= "000000";
      when 270 => pixel <= "000000";
      when 271 => pixel <= "000000";
      when 272 => pixel <= "000000";
      when 273 => pixel <= "000000";
      when 274 => pixel <= "000000";
      when 275 => pixel <= "000000";
      when 276 => pixel <= "000000";
      when 277 => pixel <= "000000";
      when 278 => pixel <= "000000";
      when 279 => pixel <= "000000";
      when 280 => pixel <= "000000";
      when 281 => pixel <= "000000";
      when 282 => pixel <= "000000";
      when 283 => pixel <= "000000";
      when 284 => pixel <= "000000";
      when 285 => pixel <= "000000";
      when 286 => pixel <= "000000";
      when 287 => pixel <= "000000";
      when 288 => pixel <= "000000";
      when 289 => pixel <= "000000";
      when 290 => pixel <= "000000";
      when 291 => pixel <= "000000";
      when 292 => pixel <= "000000";
      when 293 => pixel <= "000000";
      when 294 => pixel <= "000000";
      when 295 => pixel <= "000000";
      when 296 => pixel <= "000000";
      when 297 => pixel <= "000000";
      when 298 => pixel <= "000000";
      when 299 => pixel <= "000000";
      when 300 => pixel <= "000000";
      when 301 => pixel <= "000000";
      when 302 => pixel <= "000000";
      when 303 => pixel <= "000000";
      when 304 => pixel <= "000000";
      when 305 => pixel <= "000000";
      when 306 => pixel <= "000000";
      when 307 => pixel <= "000000";
      when 308 => pixel <= "000000";
      when 309 => pixel <= "000000";
      when 310 => pixel <= "000000";
      when 311 => pixel <= "000000";
      when 312 => pixel <= "000000";
      when 313 => pixel <= "000000";
      when 314 => pixel <= "000000";
      when 315 => pixel <= "000000";
      when 316 => pixel <= "000000";
      when 317 => pixel <= "000000";
      when 318 => pixel <= "000000";
      when 319 => pixel <= "000000";
      when 320 => pixel <= "000000";
      when 321 => pixel <= "000000";
      when 322 => pixel <= "000000";
      when 323 => pixel <= "000000";
      when 324 => pixel <= "000000";
      when 325 => pixel <= "000000";
      when 326 => pixel <= "000000";
      when 327 => pixel <= "000000";
      when 328 => pixel <= "000000";
      when 329 => pixel <= "000000";
      when 330 => pixel <= "000000";
      when 331 => pixel <= "000000";
      when 332 => pixel <= "000000";
      when 333 => pixel <= "000000";
      when 334 => pixel <= "000000";
      when 335 => pixel <= "000000";
      when 336 => pixel <= "000000";
      when 337 => pixel <= "000000";
      when 338 => pixel <= "000000";
      when 339 => pixel <= "000000";
      when 340 => pixel <= "000000";
      when 341 => pixel <= "000000";
      when 342 => pixel <= "000000";
      when 343 => pixel <= "000000";
      when 344 => pixel <= "000000";
      when 345 => pixel <= "000000";
      when 346 => pixel <= "000000";
      when 347 => pixel <= "000000";
      when 348 => pixel <= "000000";
      when 349 => pixel <= "000000";
      when 350 => pixel <= "000000";
      when 351 => pixel <= "000000";
      when 352 => pixel <= "000000";
      when 353 => pixel <= "000000";
      when 354 => pixel <= "000000";
      when 355 => pixel <= "000000";
      when 356 => pixel <= "000000";
      when 357 => pixel <= "000000";
      when 358 => pixel <= "000000";
      when 359 => pixel <= "000000";
      when 360 => pixel <= "000000";
      when 361 => pixel <= "000000";
      when 362 => pixel <= "000000";
      when 363 => pixel <= "000000";
      when 364 => pixel <= "000000";
      when 365 => pixel <= "000000";
      when 366 => pixel <= "000000";
      when 367 => pixel <= "000000";
      when 368 => pixel <= "000000";
      when 369 => pixel <= "000000";
      when 370 => pixel <= "000000";
      when 371 => pixel <= "000000";
      when 372 => pixel <= "000000";
      when 373 => pixel <= "000000";
      when 374 => pixel <= "000000";
      when 375 => pixel <= "000000";
      when 376 => pixel <= "000000";
      when 377 => pixel <= "000000";
      when 378 => pixel <= "000000";
      when 379 => pixel <= "000000";
      when 380 => pixel <= "000000";
      when 381 => pixel <= "000000";
      when 382 => pixel <= "000000";
      when 383 => pixel <= "000000";
      when 384 => pixel <= "000000";
      when 385 => pixel <= "000000";
      when 386 => pixel <= "000000";
      when 387 => pixel <= "000000";
      when 388 => pixel <= "000000";
      when 389 => pixel <= "000000";
      when 390 => pixel <= "000000";
      when 391 => pixel <= "000000";
      when 392 => pixel <= "000000";
      when 393 => pixel <= "000000";
      when 394 => pixel <= "000000";
      when 395 => pixel <= "000000";
      when 396 => pixel <= "000000";
      when 397 => pixel <= "000000";
      when 398 => pixel <= "000000";
      when 399 => pixel <= "000000";
      when 400 => pixel <= "000000";
      when 401 => pixel <= "000000";
      when 402 => pixel <= "000000";
      when 403 => pixel <= "000000";
      when 404 => pixel <= "000000";
      when 405 => pixel <= "000000";
      when 406 => pixel <= "000000";
      when 407 => pixel <= "000000";
      when 408 => pixel <= "000000";
      when 409 => pixel <= "000000";
      when 410 => pixel <= "000000";
      when 411 => pixel <= "000000";
      when 412 => pixel <= "000000";
      when 413 => pixel <= "000000";
      when 414 => pixel <= "000000";
      when 415 => pixel <= "000000";
      when 416 => pixel <= "000000";
      when 417 => pixel <= "000000";
      when 418 => pixel <= "000000";
      when 419 => pixel <= "000000";
      when 420 => pixel <= "000000";
      when 421 => pixel <= "000000";
      when 422 => pixel <= "000000";
      when 423 => pixel <= "000000";
      when 424 => pixel <= "000000";
      when 425 => pixel <= "000000";
      when 426 => pixel <= "000000";
      when 427 => pixel <= "000000";
      when 428 => pixel <= "000000";
      when 429 => pixel <= "000000";
      when 430 => pixel <= "000000";
      when 431 => pixel <= "000000";
      when 432 => pixel <= "000000";
      when 433 => pixel <= "000000";
      when 434 => pixel <= "000000";
      when 435 => pixel <= "000000";
      when 436 => pixel <= "000000";
      when 437 => pixel <= "000000";
      when 438 => pixel <= "000000";
      when 439 => pixel <= "000000";
      when 440 => pixel <= "000000";
      when 441 => pixel <= "000000";
      when 442 => pixel <= "000000";
      when 443 => pixel <= "000000";
      when 444 => pixel <= "000000";
      when 445 => pixel <= "000000";
      when 446 => pixel <= "000000";
      when 447 => pixel <= "000000";
      when 448 => pixel <= "000000";
      when 449 => pixel <= "000000";
      when 450 => pixel <= "000000";
      when 451 => pixel <= "000000";
      when 452 => pixel <= "000000";
      when 453 => pixel <= "000000";
      when 454 => pixel <= "000000";
      when 455 => pixel <= "000000";
      when 456 => pixel <= "000000";
      when 457 => pixel <= "000000";
      when 458 => pixel <= "000000";
      when 459 => pixel <= "000000";
      when 460 => pixel <= "000000";
      when 461 => pixel <= "000000";
      when 462 => pixel <= "000000";
      when 463 => pixel <= "000000";
      when 464 => pixel <= "000000";
      when 465 => pixel <= "000000";
      when 466 => pixel <= "000000";
      when 467 => pixel <= "000000";
      when 468 => pixel <= "000000";
      when 469 => pixel <= "000000";
      when 470 => pixel <= "000000";
      when 471 => pixel <= "000000";
      when 472 => pixel <= "000000";
      when 473 => pixel <= "000000";
      when 474 => pixel <= "000000";
      when 475 => pixel <= "000000";
      when 476 => pixel <= "000000";
      when 477 => pixel <= "000000";
      when 478 => pixel <= "000000";
      when 479 => pixel <= "000000";
      when 480 => pixel <= "000000";
      when 481 => pixel <= "000000";
      when 482 => pixel <= "000000";
      when 483 => pixel <= "000000";
      when 484 => pixel <= "000000";
      when 485 => pixel <= "000000";
      when 486 => pixel <= "000000";
      when 487 => pixel <= "000000";
      when 488 => pixel <= "000000";
      when 489 => pixel <= "000000";
      when 490 => pixel <= "000000";
      when 491 => pixel <= "000000";
      when 492 => pixel <= "000000";
      when 493 => pixel <= "000000";
      when 494 => pixel <= "000000";
      when 495 => pixel <= "000000";
      when 496 => pixel <= "000000";
      when 497 => pixel <= "000000";
      when 498 => pixel <= "000000";
      when 499 => pixel <= "000000";
      when 500 => pixel <= "000000";
      when 501 => pixel <= "000000";
      when 502 => pixel <= "000000";
      when 503 => pixel <= "000000";
      when 504 => pixel <= "000000";
      when 505 => pixel <= "000000";
      when 506 => pixel <= "000000";
      when 507 => pixel <= "000000";
      when 508 => pixel <= "000000";
      when 509 => pixel <= "000000";
      when 510 => pixel <= "000000";
      when 511 => pixel <= "000000";
      when 512 => pixel <= "000000";
      when 513 => pixel <= "000000";
      when 514 => pixel <= "000000";
      when 515 => pixel <= "000000";
      when 516 => pixel <= "000000";
      when 517 => pixel <= "000000";
      when 518 => pixel <= "000000";
      when 519 => pixel <= "000000";
      when 520 => pixel <= "000000";
      when 521 => pixel <= "000000";
      when 522 => pixel <= "000000";
      when 523 => pixel <= "000000";
      when 524 => pixel <= "000000";
      when 525 => pixel <= "000000";
      when 526 => pixel <= "000000";
      when 527 => pixel <= "000000";
      when 528 => pixel <= "000000";
      when 529 => pixel <= "000000";
      when 530 => pixel <= "000000";
      when 531 => pixel <= "000000";
      when 532 => pixel <= "000000";
      when 533 => pixel <= "000000";
      when 534 => pixel <= "000000";
      when 535 => pixel <= "000000";
      when 536 => pixel <= "000000";
      when 537 => pixel <= "000000";
      when 538 => pixel <= "000000";
      when 539 => pixel <= "000000";
      when 540 => pixel <= "000000";
      when 541 => pixel <= "000000";
      when 542 => pixel <= "000000";
      when 543 => pixel <= "000000";
      when 544 => pixel <= "000000";
      when 545 => pixel <= "000000";
      when 546 => pixel <= "000000";
      when 547 => pixel <= "000000";
      when 548 => pixel <= "000000";
      when 549 => pixel <= "000000";
      when 550 => pixel <= "000000";
      when 551 => pixel <= "000000";
      when 552 => pixel <= "000000";
      when 553 => pixel <= "000000";
      when 554 => pixel <= "000000";
      when 555 => pixel <= "000000";
      when 556 => pixel <= "000000";
      when 557 => pixel <= "000000";
      when 558 => pixel <= "000000";
      when 559 => pixel <= "000000";
      when 560 => pixel <= "000000";
      when 561 => pixel <= "000000";
      when 562 => pixel <= "000000";
      when 563 => pixel <= "000000";
      when 564 => pixel <= "000000";
      when 565 => pixel <= "000000";
      when 566 => pixel <= "000000";
      when 567 => pixel <= "000000";
      when 568 => pixel <= "000000";
      when 569 => pixel <= "000000";
      when 570 => pixel <= "000000";
      when 571 => pixel <= "000000";
      when 572 => pixel <= "000000";
      when 573 => pixel <= "000000";
      when 574 => pixel <= "000000";
      when 575 => pixel <= "000000";
      when 576 => pixel <= "000000";
      when 577 => pixel <= "000000";
      when 578 => pixel <= "000000";
      when 579 => pixel <= "000000";
      when 580 => pixel <= "000000";
      when 581 => pixel <= "000000";
      when 582 => pixel <= "000000";
      when 583 => pixel <= "000000";
      when 584 => pixel <= "000000";
      when 585 => pixel <= "000000";
      when 586 => pixel <= "000000";
      when 587 => pixel <= "000000";
      when 588 => pixel <= "000000";
      when 589 => pixel <= "000000";
      when 590 => pixel <= "000000";
      when 591 => pixel <= "000000";
      when 592 => pixel <= "000000";
      when 593 => pixel <= "000000";
      when 594 => pixel <= "000000";
      when 595 => pixel <= "000000";
      when 596 => pixel <= "000000";
      when 597 => pixel <= "000000";
      when 598 => pixel <= "000000";
      when 599 => pixel <= "000000";
      when 600 => pixel <= "000000";
      when 601 => pixel <= "000000";
      when 602 => pixel <= "000000";
      when 603 => pixel <= "000000";
      when 604 => pixel <= "000000";
      when 605 => pixel <= "000000";
      when 606 => pixel <= "000000";
      when 607 => pixel <= "000000";
      when 608 => pixel <= "000000";
      when 609 => pixel <= "000000";
      when 610 => pixel <= "000000";
      when 611 => pixel <= "000000";
      when 612 => pixel <= "000000";
      when 613 => pixel <= "000000";
      when 614 => pixel <= "000000";
      when 615 => pixel <= "000000";
      when 616 => pixel <= "000000";
      when 617 => pixel <= "000000";
      when 618 => pixel <= "000000";
      when 619 => pixel <= "000000";
      when 620 => pixel <= "000000";
      when 621 => pixel <= "000000";
      when 622 => pixel <= "000000";
      when 623 => pixel <= "000000";
      when 624 => pixel <= "000000";
      when 625 => pixel <= "000000";
      when 626 => pixel <= "000000";
      when 627 => pixel <= "000000";
      when 628 => pixel <= "000000";
      when 629 => pixel <= "000000";
      when 630 => pixel <= "000000";
      when 631 => pixel <= "000000";
      when 632 => pixel <= "000000";
      when 633 => pixel <= "000000";
      when 634 => pixel <= "000000";
      when 635 => pixel <= "000000";
      when 636 => pixel <= "000000";
      when 637 => pixel <= "000000";
      when 638 => pixel <= "000000";
      when 639 => pixel <= "000000";
      when 640 => pixel <= "000000";
      when 641 => pixel <= "000000";
      when 642 => pixel <= "000000";
      when 643 => pixel <= "000000";
      when 644 => pixel <= "000000";
      when 645 => pixel <= "000000";
      when 646 => pixel <= "000000";
      when 647 => pixel <= "000000";
      when 648 => pixel <= "000000";
      when 649 => pixel <= "000000";
      when 650 => pixel <= "000000";
      when 651 => pixel <= "000000";
      when 652 => pixel <= "000000";
      when 653 => pixel <= "000000";
      when 654 => pixel <= "000000";
      when 655 => pixel <= "000000";
      when 656 => pixel <= "000000";
      when 657 => pixel <= "000000";
      when 658 => pixel <= "000000";
      when 659 => pixel <= "000000";
      when 660 => pixel <= "000000";
      when 661 => pixel <= "000000";
      when 662 => pixel <= "000000";
      when 663 => pixel <= "000000";
      when 664 => pixel <= "000000";
      when 665 => pixel <= "000000";
      when 666 => pixel <= "000000";
      when 667 => pixel <= "000000";
      when 668 => pixel <= "000000";
      when 669 => pixel <= "000000";
      when 670 => pixel <= "000000";
      when 671 => pixel <= "000000";
      when 672 => pixel <= "000000";
      when 673 => pixel <= "000000";
      when 674 => pixel <= "000000";
      when 675 => pixel <= "000000";
      when 676 => pixel <= "000000";
      when 677 => pixel <= "000000";
      when 678 => pixel <= "000000";
      when 679 => pixel <= "000000";
      when 680 => pixel <= "000000";
      when 681 => pixel <= "000000";
      when 682 => pixel <= "000000";
      when 683 => pixel <= "000000";
      when 684 => pixel <= "000000";
      when 685 => pixel <= "000000";
      when 686 => pixel <= "000000";
      when 687 => pixel <= "000000";
      when 688 => pixel <= "000000";
      when 689 => pixel <= "000000";
      when 690 => pixel <= "000000";
      when 691 => pixel <= "000000";
      when 692 => pixel <= "000000";
      when 693 => pixel <= "000000";
      when 694 => pixel <= "000000";
      when 695 => pixel <= "000000";
      when 696 => pixel <= "000000";
      when 697 => pixel <= "000000";
      when 698 => pixel <= "000000";
      when 699 => pixel <= "000000";
      when 700 => pixel <= "000000";
      when 701 => pixel <= "000000";
      when 702 => pixel <= "000000";
      when 703 => pixel <= "000000";
      when 704 => pixel <= "000000";
      when 705 => pixel <= "000000";
      when 706 => pixel <= "000000";
      when 707 => pixel <= "000000";
      when 708 => pixel <= "000000";
      when 709 => pixel <= "000000";
      when 710 => pixel <= "000000";
      when 711 => pixel <= "000000";
      when 712 => pixel <= "000000";
      when 713 => pixel <= "000000";
      when 714 => pixel <= "000000";
      when 715 => pixel <= "000000";
      when 716 => pixel <= "000000";
      when 717 => pixel <= "000000";
      when 718 => pixel <= "000000";
      when 719 => pixel <= "000000";
      when 720 => pixel <= "000000";
      when 721 => pixel <= "000000";
      when 722 => pixel <= "000000";
      when 723 => pixel <= "000000";
      when 724 => pixel <= "000000";
      when 725 => pixel <= "000000";
      when 726 => pixel <= "000000";
      when 727 => pixel <= "000000";
      when 728 => pixel <= "000000";
      when 729 => pixel <= "000000";
      when 730 => pixel <= "000000";
      when 731 => pixel <= "000000";
      when 732 => pixel <= "000000";
      when 733 => pixel <= "000000";
      when 734 => pixel <= "000000";
      when 735 => pixel <= "000000";
      when 736 => pixel <= "000000";
      when 737 => pixel <= "000000";
      when 738 => pixel <= "000000";
      when 739 => pixel <= "000000";
      when 740 => pixel <= "000000";
      when 741 => pixel <= "000000";
      when 742 => pixel <= "000000";
      when 743 => pixel <= "000000";
      when 744 => pixel <= "000000";
      when 745 => pixel <= "000000";
      when 746 => pixel <= "000000";
      when 747 => pixel <= "000000";
      when 748 => pixel <= "000000";
      when 749 => pixel <= "000000";
      when 750 => pixel <= "000000";
      when 751 => pixel <= "000000";
      when 752 => pixel <= "000000";
      when 753 => pixel <= "000000";
      when 754 => pixel <= "000000";
      when 755 => pixel <= "000000";
      when 756 => pixel <= "000000";
      when 757 => pixel <= "000000";
      when 758 => pixel <= "000000";
      when 759 => pixel <= "000000";
      when 760 => pixel <= "000000";
      when 761 => pixel <= "000000";
      when 762 => pixel <= "000000";
      when 763 => pixel <= "000000";
      when 764 => pixel <= "000000";
      when 765 => pixel <= "000000";
      when 766 => pixel <= "000000";
      when 767 => pixel <= "000000";
      when 768 => pixel <= "000000";
      when 769 => pixel <= "000000";
      when 770 => pixel <= "000000";
      when 771 => pixel <= "000000";
      when 772 => pixel <= "000000";
      when 773 => pixel <= "000000";
      when 774 => pixel <= "000000";
      when 775 => pixel <= "000000";
      when 776 => pixel <= "000000";
      when 777 => pixel <= "000000";
      when 778 => pixel <= "000000";
      when 779 => pixel <= "000000";
      when 780 => pixel <= "000000";
      when 781 => pixel <= "000000";
      when 782 => pixel <= "000000";
      when 783 => pixel <= "000000";
      when 784 => pixel <= "000000";
      when 785 => pixel <= "000000";
      when 786 => pixel <= "000000";
      when 787 => pixel <= "000000";
      when 788 => pixel <= "000000";
      when 789 => pixel <= "000000";
      when 790 => pixel <= "000000";
      when 791 => pixel <= "000000";
      when 792 => pixel <= "000000";
      when 793 => pixel <= "000000";
      when 794 => pixel <= "000000";
      when 795 => pixel <= "000000";
      when 796 => pixel <= "000000";
      when 797 => pixel <= "000000";
      when 798 => pixel <= "000000";
      when 799 => pixel <= "000000";
      when 800 => pixel <= "000000";
      when 801 => pixel <= "000000";
      when 802 => pixel <= "000000";
      when 803 => pixel <= "000000";
      when 804 => pixel <= "000000";
      when 805 => pixel <= "000000";
      when 806 => pixel <= "000000";
      when 807 => pixel <= "000000";
      when 808 => pixel <= "000000";
      when 809 => pixel <= "000000";
      when 810 => pixel <= "000000";
      when 811 => pixel <= "000000";
      when 812 => pixel <= "000000";
      when 813 => pixel <= "000000";
      when 814 => pixel <= "000000";
      when 815 => pixel <= "000000";
      when 816 => pixel <= "000000";
      when 817 => pixel <= "000000";
      when 818 => pixel <= "000000";
      when 819 => pixel <= "000000";
      when 820 => pixel <= "000000";
      when 821 => pixel <= "000000";
      when 822 => pixel <= "000000";
      when 823 => pixel <= "000000";
      when 824 => pixel <= "000000";
      when 825 => pixel <= "000000";
      when 826 => pixel <= "000000";
      when 827 => pixel <= "000000";
      when 828 => pixel <= "000000";
      when 829 => pixel <= "000000";
      when 830 => pixel <= "000000";
      when 831 => pixel <= "000000";
      when 832 => pixel <= "000000";
      when 833 => pixel <= "000000";
      when 834 => pixel <= "000000";
      when 835 => pixel <= "000000";
      when 836 => pixel <= "000000";
      when 837 => pixel <= "000000";
      when 838 => pixel <= "000000";
      when 839 => pixel <= "000000";
      when 840 => pixel <= "000000";
      when 841 => pixel <= "000000";
      when 842 => pixel <= "000000";
      when 843 => pixel <= "000000";
      when 844 => pixel <= "000000";
      when 845 => pixel <= "000000";
      when 846 => pixel <= "000000";
      when 847 => pixel <= "000000";
      when 848 => pixel <= "000000";
      when 849 => pixel <= "000000";
      when 850 => pixel <= "000000";
      when 851 => pixel <= "000000";
      when 852 => pixel <= "000000";
      when 853 => pixel <= "000000";
      when 854 => pixel <= "000000";
      when 855 => pixel <= "000000";
      when 856 => pixel <= "000000";
      when 857 => pixel <= "000000";
      when 858 => pixel <= "000000";
      when 859 => pixel <= "000000";
      when 860 => pixel <= "000000";
      when 861 => pixel <= "000000";
      when 862 => pixel <= "000000";
      when 863 => pixel <= "000000";
      when 864 => pixel <= "000000";
      when 865 => pixel <= "000000";
      when 866 => pixel <= "000000";
      when 867 => pixel <= "000000";
      when 868 => pixel <= "000000";
      when 869 => pixel <= "000000";
      when 870 => pixel <= "000000";
      when 871 => pixel <= "000000";
      when 872 => pixel <= "000000";
      when 873 => pixel <= "000000";
      when 874 => pixel <= "000000";
      when 875 => pixel <= "000000";
      when 876 => pixel <= "000000";
      when 877 => pixel <= "000000";
      when 878 => pixel <= "000000";
      when 879 => pixel <= "000000";
      when 880 => pixel <= "000000";
      when 881 => pixel <= "000000";
      when 882 => pixel <= "000000";
      when 883 => pixel <= "000000";
      when 884 => pixel <= "000000";
      when 885 => pixel <= "000000";
      when 886 => pixel <= "000000";
      when 887 => pixel <= "000000";
      when 888 => pixel <= "000000";
      when 889 => pixel <= "000000";
      when 890 => pixel <= "000000";
      when 891 => pixel <= "000000";
      when 892 => pixel <= "000000";
      when 893 => pixel <= "000000";
      when 894 => pixel <= "000000";
      when 895 => pixel <= "000000";
      when 896 => pixel <= "000000";
      when 897 => pixel <= "000000";
      when 898 => pixel <= "000000";
      when 899 => pixel <= "000000";
      when 900 => pixel <= "000000";
      when 901 => pixel <= "000000";
      when 902 => pixel <= "000000";
      when 903 => pixel <= "000000";
      when 904 => pixel <= "000000";
      when 905 => pixel <= "000000";
      when 906 => pixel <= "000000";
      when 907 => pixel <= "000000";
      when 908 => pixel <= "000000";
      when 909 => pixel <= "000000";
      when 910 => pixel <= "000000";
      when 911 => pixel <= "000000";
      when 912 => pixel <= "000000";
      when 913 => pixel <= "000000";
      when 914 => pixel <= "000000";
      when 915 => pixel <= "000000";
      when 916 => pixel <= "000000";
      when 917 => pixel <= "000000";
      when 918 => pixel <= "000000";
      when 919 => pixel <= "000000";
      when 920 => pixel <= "000000";
      when 921 => pixel <= "000000";
      when 922 => pixel <= "000000";
      when 923 => pixel <= "000000";
      when 924 => pixel <= "000000";
      when 925 => pixel <= "000000";
      when 926 => pixel <= "000000";
      when 927 => pixel <= "000000";
      when 928 => pixel <= "000000";
      when 929 => pixel <= "000000";
      when 930 => pixel <= "000000";
      when 931 => pixel <= "000000";
      when 932 => pixel <= "000000";
      when 933 => pixel <= "000000";
      when 934 => pixel <= "000000";
      when 935 => pixel <= "000000";
      when 936 => pixel <= "000000";
      when 937 => pixel <= "000000";
      when 938 => pixel <= "000000";
      when 939 => pixel <= "000000";
      when 940 => pixel <= "000000";
      when 941 => pixel <= "000000";
      when 942 => pixel <= "000000";
      when 943 => pixel <= "000000";
      when 944 => pixel <= "000000";
      when 945 => pixel <= "000000";
      when 946 => pixel <= "000000";
      when 947 => pixel <= "000000";
      when 948 => pixel <= "000000";
      when 949 => pixel <= "000000";
      when 950 => pixel <= "000000";
      when 951 => pixel <= "000000";
      when 952 => pixel <= "000000";
      when 953 => pixel <= "000000";
      when 954 => pixel <= "000000";
      when 955 => pixel <= "000000";
      when 956 => pixel <= "000000";
      when 957 => pixel <= "000000";
      when 958 => pixel <= "000000";
      when 959 => pixel <= "000000";
      when 960 => pixel <= "000000";
      when 961 => pixel <= "000000";
      when 962 => pixel <= "000000";
      when 963 => pixel <= "000000";
      when 964 => pixel <= "000000";
      when 965 => pixel <= "000000";
      when 966 => pixel <= "000000";
      when 967 => pixel <= "000000";
      when 968 => pixel <= "000000";
      when 969 => pixel <= "000000";
      when 970 => pixel <= "000000";
      when 971 => pixel <= "000000";
      when 972 => pixel <= "000000";
      when 973 => pixel <= "000000";
      when 974 => pixel <= "000000";
      when 975 => pixel <= "000000";
      when 976 => pixel <= "000000";
      when 977 => pixel <= "000000";
      when 978 => pixel <= "000000";
      when 979 => pixel <= "000000";
      when 980 => pixel <= "000000";
      when 981 => pixel <= "000000";
      when 982 => pixel <= "000000";
      when 983 => pixel <= "000000";
      when 984 => pixel <= "000000";
      when 985 => pixel <= "000000";
      when 986 => pixel <= "000000";
      when 987 => pixel <= "000000";
      when 988 => pixel <= "000000";
      when 989 => pixel <= "000000";
      when 990 => pixel <= "000000";
      when 991 => pixel <= "000000";
      when 992 => pixel <= "000000";
      when 993 => pixel <= "000000";
      when 994 => pixel <= "000000";
      when 995 => pixel <= "000000";
      when 996 => pixel <= "000000";
      when 997 => pixel <= "000000";
      when 998 => pixel <= "000000";
      when 999 => pixel <= "000000";
      when 1000 => pixel <= "000000";
      when 1001 => pixel <= "000000";
      when 1002 => pixel <= "000000";
      when 1003 => pixel <= "000000";
      when 1004 => pixel <= "000000";
      when 1005 => pixel <= "000000";
      when 1006 => pixel <= "000000";
      when 1007 => pixel <= "000000";
      when 1008 => pixel <= "000000";
      when 1009 => pixel <= "000000";
      when 1010 => pixel <= "000000";
      when 1011 => pixel <= "000000";
      when 1012 => pixel <= "000000";
      when 1013 => pixel <= "000000";
      when 1014 => pixel <= "000000";
      when 1015 => pixel <= "000000";
      when 1016 => pixel <= "000000";
      when 1017 => pixel <= "000000";
      when 1018 => pixel <= "000000";
      when 1019 => pixel <= "000000";
      when 1020 => pixel <= "000000";
      when 1021 => pixel <= "000000";
      when 1022 => pixel <= "000000";
      when 1023 => pixel <= "000000";
      when 1024 => pixel <= "000000";
      when 1025 => pixel <= "000000";
      when 1026 => pixel <= "000000";
      when 1027 => pixel <= "000000";
      when 1028 => pixel <= "000000";
      when 1029 => pixel <= "000000";
      when 1030 => pixel <= "000000";
      when 1031 => pixel <= "000000";
      when 1032 => pixel <= "000000";
      when 1033 => pixel <= "000000";
      when 1034 => pixel <= "000000";
      when 1035 => pixel <= "000000";
      when 1036 => pixel <= "000000";
      when 1037 => pixel <= "000000";
      when 1038 => pixel <= "000000";
      when 1039 => pixel <= "000000";
      when 1040 => pixel <= "000000";
      when 1041 => pixel <= "000000";
      when 1042 => pixel <= "000000";
      when 1043 => pixel <= "000000";
      when 1044 => pixel <= "000000";
      when 1045 => pixel <= "000000";
      when 1046 => pixel <= "000000";
      when 1047 => pixel <= "000000";
      when 1048 => pixel <= "000000";
      when 1049 => pixel <= "000000";
      when 1050 => pixel <= "000000";
      when 1051 => pixel <= "000000";
      when 1052 => pixel <= "000000";
      when 1053 => pixel <= "000000";
      when 1054 => pixel <= "000000";
      when 1055 => pixel <= "000000";
      when 1056 => pixel <= "000000";
      when 1057 => pixel <= "000000";
      when 1058 => pixel <= "000000";
      when 1059 => pixel <= "000000";
      when 1060 => pixel <= "000000";
      when 1061 => pixel <= "000000";
      when 1062 => pixel <= "000000";
      when 1063 => pixel <= "000000";
      when 1064 => pixel <= "000000";
      when 1065 => pixel <= "000000";
      when 1066 => pixel <= "000000";
      when 1067 => pixel <= "000000";
      when 1068 => pixel <= "000000";
      when 1069 => pixel <= "000000";
      when 1070 => pixel <= "000000";
      when 1071 => pixel <= "000000";
      when 1072 => pixel <= "000000";
      when 1073 => pixel <= "000000";
      when 1074 => pixel <= "000000";
      when 1075 => pixel <= "000000";
      when 1076 => pixel <= "000000";
      when 1077 => pixel <= "000000";
      when 1078 => pixel <= "000000";
      when 1079 => pixel <= "000000";
      when 1080 => pixel <= "000000";
      when 1081 => pixel <= "000000";
      when 1082 => pixel <= "000000";
      when 1083 => pixel <= "000000";
      when 1084 => pixel <= "000000";
      when 1085 => pixel <= "000000";
      when 1086 => pixel <= "000000";
      when 1087 => pixel <= "000000";
      when 1088 => pixel <= "000000";
      when 1089 => pixel <= "000000";
      when 1090 => pixel <= "000000";
      when 1091 => pixel <= "000000";
      when 1092 => pixel <= "000000";
      when 1093 => pixel <= "000000";
      when 1094 => pixel <= "000000";
      when 1095 => pixel <= "000000";
      when 1096 => pixel <= "000000";
      when 1097 => pixel <= "000000";
      when 1098 => pixel <= "000000";
      when 1099 => pixel <= "000000";
      when 1100 => pixel <= "000000";
      when 1101 => pixel <= "000000";
      when 1102 => pixel <= "000000";
      when 1103 => pixel <= "000000";
      when 1104 => pixel <= "000000";
      when 1105 => pixel <= "000000";
      when 1106 => pixel <= "000000";
      when 1107 => pixel <= "000000";
      when 1108 => pixel <= "000000";
      when 1109 => pixel <= "000000";
      when 1110 => pixel <= "000000";
      when 1111 => pixel <= "000000";
      when 1112 => pixel <= "000000";
      when 1113 => pixel <= "000000";
      when 1114 => pixel <= "000000";
      when 1115 => pixel <= "000000";
      when 1116 => pixel <= "000000";
      when 1117 => pixel <= "000000";
      when 1118 => pixel <= "000000";
      when 1119 => pixel <= "000000";
      when 1120 => pixel <= "000000";
      when 1121 => pixel <= "000000";
      when 1122 => pixel <= "000000";
      when 1123 => pixel <= "000000";
      when 1124 => pixel <= "000000";
      when 1125 => pixel <= "000000";
      when 1126 => pixel <= "000000";
      when 1127 => pixel <= "000000";
      when 1128 => pixel <= "000000";
      when 1129 => pixel <= "000000";
      when 1130 => pixel <= "000000";
      when 1131 => pixel <= "000000";
      when 1132 => pixel <= "000000";
      when 1133 => pixel <= "000000";
      when 1134 => pixel <= "000000";
      when 1135 => pixel <= "000000";
      when 1136 => pixel <= "000000";
      when 1137 => pixel <= "000000";
      when 1138 => pixel <= "000000";
      when 1139 => pixel <= "000000";
      when 1140 => pixel <= "000000";
      when 1141 => pixel <= "000000";
      when 1142 => pixel <= "000000";
      when 1143 => pixel <= "000000";
      when 1144 => pixel <= "000000";
      when 1145 => pixel <= "000000";
      when 1146 => pixel <= "000000";
      when 1147 => pixel <= "000000";
      when 1148 => pixel <= "000000";
      when 1149 => pixel <= "000000";
      when 1150 => pixel <= "000000";
      when 1151 => pixel <= "000000";
      when 1152 => pixel <= "000000";
      when 1153 => pixel <= "000000";
      when 1154 => pixel <= "000000";
      when 1155 => pixel <= "000000";
      when 1156 => pixel <= "001101";
      when 1157 => pixel <= "001101";
      when 1158 => pixel <= "001101";
      when 1159 => pixel <= "001101";
      when 1160 => pixel <= "000000";
      when 1161 => pixel <= "000000";
      when 1162 => pixel <= "000000";
      when 1163 => pixel <= "000000";
      when 1164 => pixel <= "000000";
      when 1165 => pixel <= "000000";
      when 1166 => pixel <= "001101";
      when 1167 => pixel <= "000000";
      when 1168 => pixel <= "000000";
      when 1169 => pixel <= "000000";
      when 1170 => pixel <= "000000";
      when 1171 => pixel <= "000000";
      when 1172 => pixel <= "001101";
      when 1173 => pixel <= "001101";
      when 1174 => pixel <= "000000";
      when 1175 => pixel <= "000000";
      when 1176 => pixel <= "000000";
      when 1177 => pixel <= "001101";
      when 1178 => pixel <= "001101";
      when 1179 => pixel <= "000000";
      when 1180 => pixel <= "000000";
      when 1181 => pixel <= "001101";
      when 1182 => pixel <= "001101";
      when 1183 => pixel <= "001101";
      when 1184 => pixel <= "001101";
      when 1185 => pixel <= "001101";
      when 1186 => pixel <= "001101";
      when 1187 => pixel <= "001101";
      when 1188 => pixel <= "000000";
      when 1189 => pixel <= "000000";
      when 1190 => pixel <= "000000";
      when 1191 => pixel <= "000000";
      when 1192 => pixel <= "000000";
      when 1193 => pixel <= "000000";
      when 1194 => pixel <= "000000";
      when 1195 => pixel <= "000000";
      when 1196 => pixel <= "000000";
      when 1197 => pixel <= "000000";
      when 1198 => pixel <= "000000";
      when 1199 => pixel <= "000000";
      when 1200 => pixel <= "000000";
      when 1201 => pixel <= "001101";
      when 1202 => pixel <= "001101";
      when 1203 => pixel <= "001101";
      when 1204 => pixel <= "001101";
      when 1205 => pixel <= "001101";
      when 1206 => pixel <= "000000";
      when 1207 => pixel <= "000000";
      when 1208 => pixel <= "000000";
      when 1209 => pixel <= "001101";
      when 1210 => pixel <= "001101";
      when 1211 => pixel <= "000000";
      when 1212 => pixel <= "000000";
      when 1213 => pixel <= "000000";
      when 1214 => pixel <= "001101";
      when 1215 => pixel <= "001101";
      when 1216 => pixel <= "000000";
      when 1217 => pixel <= "000000";
      when 1218 => pixel <= "001101";
      when 1219 => pixel <= "001101";
      when 1220 => pixel <= "001101";
      when 1221 => pixel <= "001101";
      when 1222 => pixel <= "001101";
      when 1223 => pixel <= "001101";
      when 1224 => pixel <= "001101";
      when 1225 => pixel <= "000000";
      when 1226 => pixel <= "000000";
      when 1227 => pixel <= "001101";
      when 1228 => pixel <= "001101";
      when 1229 => pixel <= "001101";
      when 1230 => pixel <= "001101";
      when 1231 => pixel <= "001101";
      when 1232 => pixel <= "001101";
      when 1233 => pixel <= "000000";
      when 1234 => pixel <= "000000";
      when 1235 => pixel <= "000000";
      when 1236 => pixel <= "000000";
      when 1237 => pixel <= "000000";
      when 1238 => pixel <= "000000";
      when 1239 => pixel <= "001101";
      when 1240 => pixel <= "001101";
      when 1241 => pixel <= "000000";
      when 1242 => pixel <= "000000";
      when 1243 => pixel <= "000000";
      when 1244 => pixel <= "000000";
      when 1245 => pixel <= "000000";
      when 1246 => pixel <= "000000";
      when 1247 => pixel <= "000000";
      when 1248 => pixel <= "000000";
      when 1249 => pixel <= "000000";
      when 1250 => pixel <= "000000";
      when 1251 => pixel <= "000000";
      when 1252 => pixel <= "000000";
      when 1253 => pixel <= "000000";
      when 1254 => pixel <= "000000";
      when 1255 => pixel <= "000000";
      when 1256 => pixel <= "000000";
      when 1257 => pixel <= "000000";
      when 1258 => pixel <= "000000";
      when 1259 => pixel <= "000000";
      when 1260 => pixel <= "000000";
      when 1261 => pixel <= "000000";
      when 1262 => pixel <= "000000";
      when 1263 => pixel <= "000000";
      when 1264 => pixel <= "000000";
      when 1265 => pixel <= "000000";
      when 1266 => pixel <= "000000";
      when 1267 => pixel <= "000000";
      when 1268 => pixel <= "000000";
      when 1269 => pixel <= "000000";
      when 1270 => pixel <= "000000";
      when 1271 => pixel <= "000000";
      when 1272 => pixel <= "000000";
      when 1273 => pixel <= "000000";
      when 1274 => pixel <= "000000";
      when 1275 => pixel <= "000000";
      when 1276 => pixel <= "000000";
      when 1277 => pixel <= "000000";
      when 1278 => pixel <= "000000";
      when 1279 => pixel <= "000000";
      when 1280 => pixel <= "000000";
      when 1281 => pixel <= "000000";
      when 1282 => pixel <= "000000";
      when 1283 => pixel <= "000000";
      when 1284 => pixel <= "000000";
      when 1285 => pixel <= "000000";
      when 1286 => pixel <= "000000";
      when 1287 => pixel <= "000000";
      when 1288 => pixel <= "000000";
      when 1289 => pixel <= "000000";
      when 1290 => pixel <= "000000";
      when 1291 => pixel <= "000000";
      when 1292 => pixel <= "000000";
      when 1293 => pixel <= "000000";
      when 1294 => pixel <= "000000";
      when 1295 => pixel <= "000000";
      when 1296 => pixel <= "000000";
      when 1297 => pixel <= "000000";
      when 1298 => pixel <= "000000";
      when 1299 => pixel <= "000000";
      when 1300 => pixel <= "000000";
      when 1301 => pixel <= "000000";
      when 1302 => pixel <= "000000";
      when 1303 => pixel <= "000000";
      when 1304 => pixel <= "000000";
      when 1305 => pixel <= "000000";
      when 1306 => pixel <= "000000";
      when 1307 => pixel <= "000000";
      when 1308 => pixel <= "000000";
      when 1309 => pixel <= "000000";
      when 1310 => pixel <= "000000";
      when 1311 => pixel <= "000000";
      when 1312 => pixel <= "000000";
      when 1313 => pixel <= "000000";
      when 1314 => pixel <= "000000";
      when 1315 => pixel <= "001101";
      when 1316 => pixel <= "001101";
      when 1317 => pixel <= "000000";
      when 1318 => pixel <= "000000";
      when 1319 => pixel <= "001101";
      when 1320 => pixel <= "001101";
      when 1321 => pixel <= "000000";
      when 1322 => pixel <= "000000";
      when 1323 => pixel <= "000000";
      when 1324 => pixel <= "000000";
      when 1325 => pixel <= "001101";
      when 1326 => pixel <= "001101";
      when 1327 => pixel <= "001101";
      when 1328 => pixel <= "000000";
      when 1329 => pixel <= "000000";
      when 1330 => pixel <= "000000";
      when 1331 => pixel <= "000000";
      when 1332 => pixel <= "001101";
      when 1333 => pixel <= "001101";
      when 1334 => pixel <= "001101";
      when 1335 => pixel <= "000000";
      when 1336 => pixel <= "001101";
      when 1337 => pixel <= "001101";
      when 1338 => pixel <= "001101";
      when 1339 => pixel <= "000000";
      when 1340 => pixel <= "000000";
      when 1341 => pixel <= "000000";
      when 1342 => pixel <= "001101";
      when 1343 => pixel <= "001101";
      when 1344 => pixel <= "000000";
      when 1345 => pixel <= "000000";
      when 1346 => pixel <= "001101";
      when 1347 => pixel <= "001101";
      when 1348 => pixel <= "000000";
      when 1349 => pixel <= "000000";
      when 1350 => pixel <= "000000";
      when 1351 => pixel <= "000000";
      when 1352 => pixel <= "000000";
      when 1353 => pixel <= "000000";
      when 1354 => pixel <= "000000";
      when 1355 => pixel <= "000000";
      when 1356 => pixel <= "000000";
      when 1357 => pixel <= "000000";
      when 1358 => pixel <= "000000";
      when 1359 => pixel <= "001101";
      when 1360 => pixel <= "001101";
      when 1361 => pixel <= "001101";
      when 1362 => pixel <= "000000";
      when 1363 => pixel <= "000000";
      when 1364 => pixel <= "000000";
      when 1365 => pixel <= "001101";
      when 1366 => pixel <= "001101";
      when 1367 => pixel <= "000000";
      when 1368 => pixel <= "000000";
      when 1369 => pixel <= "001101";
      when 1370 => pixel <= "001101";
      when 1371 => pixel <= "000000";
      when 1372 => pixel <= "000000";
      when 1373 => pixel <= "000000";
      when 1374 => pixel <= "001101";
      when 1375 => pixel <= "001101";
      when 1376 => pixel <= "000000";
      when 1377 => pixel <= "000000";
      when 1378 => pixel <= "000000";
      when 1379 => pixel <= "001101";
      when 1380 => pixel <= "001101";
      when 1381 => pixel <= "000000";
      when 1382 => pixel <= "000000";
      when 1383 => pixel <= "001101";
      when 1384 => pixel <= "001101";
      when 1385 => pixel <= "000000";
      when 1386 => pixel <= "000000";
      when 1387 => pixel <= "000000";
      when 1388 => pixel <= "001101";
      when 1389 => pixel <= "001101";
      when 1390 => pixel <= "000000";
      when 1391 => pixel <= "000000";
      when 1392 => pixel <= "001101";
      when 1393 => pixel <= "001101";
      when 1394 => pixel <= "000000";
      when 1395 => pixel <= "000000";
      when 1396 => pixel <= "000000";
      when 1397 => pixel <= "000000";
      when 1398 => pixel <= "001101";
      when 1399 => pixel <= "001101";
      when 1400 => pixel <= "001101";
      when 1401 => pixel <= "001101";
      when 1402 => pixel <= "000000";
      when 1403 => pixel <= "000000";
      when 1404 => pixel <= "000000";
      when 1405 => pixel <= "000000";
      when 1406 => pixel <= "000000";
      when 1407 => pixel <= "000000";
      when 1408 => pixel <= "000000";
      when 1409 => pixel <= "000000";
      when 1410 => pixel <= "000000";
      when 1411 => pixel <= "000000";
      when 1412 => pixel <= "000000";
      when 1413 => pixel <= "000000";
      when 1414 => pixel <= "000000";
      when 1415 => pixel <= "000000";
      when 1416 => pixel <= "000000";
      when 1417 => pixel <= "000000";
      when 1418 => pixel <= "000000";
      when 1419 => pixel <= "000000";
      when 1420 => pixel <= "000000";
      when 1421 => pixel <= "000000";
      when 1422 => pixel <= "000000";
      when 1423 => pixel <= "000000";
      when 1424 => pixel <= "000000";
      when 1425 => pixel <= "000000";
      when 1426 => pixel <= "000000";
      when 1427 => pixel <= "000000";
      when 1428 => pixel <= "000000";
      when 1429 => pixel <= "000000";
      when 1430 => pixel <= "000000";
      when 1431 => pixel <= "000000";
      when 1432 => pixel <= "000000";
      when 1433 => pixel <= "000000";
      when 1434 => pixel <= "000000";
      when 1435 => pixel <= "000000";
      when 1436 => pixel <= "000000";
      when 1437 => pixel <= "000000";
      when 1438 => pixel <= "000000";
      when 1439 => pixel <= "000000";
      when 1440 => pixel <= "000000";
      when 1441 => pixel <= "000000";
      when 1442 => pixel <= "000000";
      when 1443 => pixel <= "000000";
      when 1444 => pixel <= "000000";
      when 1445 => pixel <= "000000";
      when 1446 => pixel <= "000000";
      when 1447 => pixel <= "000000";
      when 1448 => pixel <= "000000";
      when 1449 => pixel <= "000000";
      when 1450 => pixel <= "000000";
      when 1451 => pixel <= "000000";
      when 1452 => pixel <= "000000";
      when 1453 => pixel <= "000000";
      when 1454 => pixel <= "000000";
      when 1455 => pixel <= "000000";
      when 1456 => pixel <= "000000";
      when 1457 => pixel <= "000000";
      when 1458 => pixel <= "000000";
      when 1459 => pixel <= "000000";
      when 1460 => pixel <= "000000";
      when 1461 => pixel <= "000000";
      when 1462 => pixel <= "000000";
      when 1463 => pixel <= "000000";
      when 1464 => pixel <= "000000";
      when 1465 => pixel <= "000000";
      when 1466 => pixel <= "000000";
      when 1467 => pixel <= "000000";
      when 1468 => pixel <= "000000";
      when 1469 => pixel <= "000000";
      when 1470 => pixel <= "000000";
      when 1471 => pixel <= "000000";
      when 1472 => pixel <= "000000";
      when 1473 => pixel <= "000000";
      when 1474 => pixel <= "001101";
      when 1475 => pixel <= "001101";
      when 1476 => pixel <= "000000";
      when 1477 => pixel <= "000000";
      when 1478 => pixel <= "000000";
      when 1479 => pixel <= "000000";
      when 1480 => pixel <= "001101";
      when 1481 => pixel <= "000000";
      when 1482 => pixel <= "000000";
      when 1483 => pixel <= "000000";
      when 1484 => pixel <= "001101";
      when 1485 => pixel <= "001101";
      when 1486 => pixel <= "000000";
      when 1487 => pixel <= "001101";
      when 1488 => pixel <= "001101";
      when 1489 => pixel <= "000000";
      when 1490 => pixel <= "000000";
      when 1491 => pixel <= "000000";
      when 1492 => pixel <= "001101";
      when 1493 => pixel <= "001101";
      when 1494 => pixel <= "001101";
      when 1495 => pixel <= "001101";
      when 1496 => pixel <= "001101";
      when 1497 => pixel <= "001101";
      when 1498 => pixel <= "001101";
      when 1499 => pixel <= "000000";
      when 1500 => pixel <= "000000";
      when 1501 => pixel <= "000000";
      when 1502 => pixel <= "001101";
      when 1503 => pixel <= "001101";
      when 1504 => pixel <= "000000";
      when 1505 => pixel <= "000000";
      when 1506 => pixel <= "000000";
      when 1507 => pixel <= "001101";
      when 1508 => pixel <= "000000";
      when 1509 => pixel <= "000000";
      when 1510 => pixel <= "000000";
      when 1511 => pixel <= "000000";
      when 1512 => pixel <= "000000";
      when 1513 => pixel <= "000000";
      when 1514 => pixel <= "000000";
      when 1515 => pixel <= "000000";
      when 1516 => pixel <= "000000";
      when 1517 => pixel <= "000000";
      when 1518 => pixel <= "000000";
      when 1519 => pixel <= "001101";
      when 1520 => pixel <= "001101";
      when 1521 => pixel <= "001101";
      when 1522 => pixel <= "000000";
      when 1523 => pixel <= "000000";
      when 1524 => pixel <= "000000";
      when 1525 => pixel <= "001101";
      when 1526 => pixel <= "001101";
      when 1527 => pixel <= "000000";
      when 1528 => pixel <= "000000";
      when 1529 => pixel <= "001101";
      when 1530 => pixel <= "001101";
      when 1531 => pixel <= "000000";
      when 1532 => pixel <= "000000";
      when 1533 => pixel <= "000000";
      when 1534 => pixel <= "001101";
      when 1535 => pixel <= "001101";
      when 1536 => pixel <= "000000";
      when 1537 => pixel <= "000000";
      when 1538 => pixel <= "000000";
      when 1539 => pixel <= "001101";
      when 1540 => pixel <= "001101";
      when 1541 => pixel <= "000000";
      when 1542 => pixel <= "000000";
      when 1543 => pixel <= "000000";
      when 1544 => pixel <= "001101";
      when 1545 => pixel <= "000000";
      when 1546 => pixel <= "000000";
      when 1547 => pixel <= "000000";
      when 1548 => pixel <= "001101";
      when 1549 => pixel <= "001101";
      when 1550 => pixel <= "000000";
      when 1551 => pixel <= "000000";
      when 1552 => pixel <= "001101";
      when 1553 => pixel <= "001101";
      when 1554 => pixel <= "000000";
      when 1555 => pixel <= "000000";
      when 1556 => pixel <= "000000";
      when 1557 => pixel <= "000000";
      when 1558 => pixel <= "001101";
      when 1559 => pixel <= "001101";
      when 1560 => pixel <= "001101";
      when 1561 => pixel <= "001101";
      when 1562 => pixel <= "000000";
      when 1563 => pixel <= "000000";
      when 1564 => pixel <= "000000";
      when 1565 => pixel <= "000000";
      when 1566 => pixel <= "000000";
      when 1567 => pixel <= "000000";
      when 1568 => pixel <= "000000";
      when 1569 => pixel <= "000000";
      when 1570 => pixel <= "000000";
      when 1571 => pixel <= "000000";
      when 1572 => pixel <= "000000";
      when 1573 => pixel <= "000000";
      when 1574 => pixel <= "000000";
      when 1575 => pixel <= "000000";
      when 1576 => pixel <= "000000";
      when 1577 => pixel <= "000000";
      when 1578 => pixel <= "000000";
      when 1579 => pixel <= "000000";
      when 1580 => pixel <= "000000";
      when 1581 => pixel <= "000000";
      when 1582 => pixel <= "000000";
      when 1583 => pixel <= "000000";
      when 1584 => pixel <= "000000";
      when 1585 => pixel <= "000000";
      when 1586 => pixel <= "000000";
      when 1587 => pixel <= "000000";
      when 1588 => pixel <= "000000";
      when 1589 => pixel <= "000000";
      when 1590 => pixel <= "000000";
      when 1591 => pixel <= "000000";
      when 1592 => pixel <= "000000";
      when 1593 => pixel <= "000000";
      when 1594 => pixel <= "000000";
      when 1595 => pixel <= "000000";
      when 1596 => pixel <= "000000";
      when 1597 => pixel <= "000000";
      when 1598 => pixel <= "000000";
      when 1599 => pixel <= "000000";
      when 1600 => pixel <= "000000";
      when 1601 => pixel <= "000000";
      when 1602 => pixel <= "000000";
      when 1603 => pixel <= "000000";
      when 1604 => pixel <= "000000";
      when 1605 => pixel <= "000000";
      when 1606 => pixel <= "000000";
      when 1607 => pixel <= "000000";
      when 1608 => pixel <= "000000";
      when 1609 => pixel <= "000000";
      when 1610 => pixel <= "000000";
      when 1611 => pixel <= "000000";
      when 1612 => pixel <= "000000";
      when 1613 => pixel <= "000000";
      when 1614 => pixel <= "000000";
      when 1615 => pixel <= "000000";
      when 1616 => pixel <= "000000";
      when 1617 => pixel <= "000000";
      when 1618 => pixel <= "000000";
      when 1619 => pixel <= "000000";
      when 1620 => pixel <= "000000";
      when 1621 => pixel <= "000000";
      when 1622 => pixel <= "000000";
      when 1623 => pixel <= "000000";
      when 1624 => pixel <= "000000";
      when 1625 => pixel <= "000000";
      when 1626 => pixel <= "000000";
      when 1627 => pixel <= "000000";
      when 1628 => pixel <= "000000";
      when 1629 => pixel <= "000000";
      when 1630 => pixel <= "000000";
      when 1631 => pixel <= "000000";
      when 1632 => pixel <= "000000";
      when 1633 => pixel <= "000000";
      when 1634 => pixel <= "001101";
      when 1635 => pixel <= "001101";
      when 1636 => pixel <= "000000";
      when 1637 => pixel <= "000000";
      when 1638 => pixel <= "000000";
      when 1639 => pixel <= "000000";
      when 1640 => pixel <= "000000";
      when 1641 => pixel <= "000000";
      when 1642 => pixel <= "000000";
      when 1643 => pixel <= "001101";
      when 1644 => pixel <= "001101";
      when 1645 => pixel <= "000000";
      when 1646 => pixel <= "000000";
      when 1647 => pixel <= "000000";
      when 1648 => pixel <= "001101";
      when 1649 => pixel <= "001101";
      when 1650 => pixel <= "000000";
      when 1651 => pixel <= "000000";
      when 1652 => pixel <= "001101";
      when 1653 => pixel <= "001101";
      when 1654 => pixel <= "001101";
      when 1655 => pixel <= "001101";
      when 1656 => pixel <= "001101";
      when 1657 => pixel <= "001101";
      when 1658 => pixel <= "001101";
      when 1659 => pixel <= "000000";
      when 1660 => pixel <= "000000";
      when 1661 => pixel <= "000000";
      when 1662 => pixel <= "001101";
      when 1663 => pixel <= "001101";
      when 1664 => pixel <= "000000";
      when 1665 => pixel <= "001101";
      when 1666 => pixel <= "000000";
      when 1667 => pixel <= "000000";
      when 1668 => pixel <= "000000";
      when 1669 => pixel <= "000000";
      when 1670 => pixel <= "000000";
      when 1671 => pixel <= "000000";
      when 1672 => pixel <= "000000";
      when 1673 => pixel <= "000000";
      when 1674 => pixel <= "000000";
      when 1675 => pixel <= "000000";
      when 1676 => pixel <= "000000";
      when 1677 => pixel <= "000000";
      when 1678 => pixel <= "000000";
      when 1679 => pixel <= "001101";
      when 1680 => pixel <= "001101";
      when 1681 => pixel <= "001101";
      when 1682 => pixel <= "000000";
      when 1683 => pixel <= "000000";
      when 1684 => pixel <= "000000";
      when 1685 => pixel <= "001101";
      when 1686 => pixel <= "001101";
      when 1687 => pixel <= "000000";
      when 1688 => pixel <= "000000";
      when 1689 => pixel <= "001101";
      when 1690 => pixel <= "001101";
      when 1691 => pixel <= "000000";
      when 1692 => pixel <= "000000";
      when 1693 => pixel <= "000000";
      when 1694 => pixel <= "001101";
      when 1695 => pixel <= "001101";
      when 1696 => pixel <= "000000";
      when 1697 => pixel <= "000000";
      when 1698 => pixel <= "000000";
      when 1699 => pixel <= "001101";
      when 1700 => pixel <= "001101";
      when 1701 => pixel <= "000000";
      when 1702 => pixel <= "001101";
      when 1703 => pixel <= "000000";
      when 1704 => pixel <= "000000";
      when 1705 => pixel <= "000000";
      when 1706 => pixel <= "000000";
      when 1707 => pixel <= "000000";
      when 1708 => pixel <= "001101";
      when 1709 => pixel <= "001101";
      when 1710 => pixel <= "000000";
      when 1711 => pixel <= "000000";
      when 1712 => pixel <= "001101";
      when 1713 => pixel <= "001101";
      when 1714 => pixel <= "000000";
      when 1715 => pixel <= "000000";
      when 1716 => pixel <= "000000";
      when 1717 => pixel <= "000000";
      when 1718 => pixel <= "001101";
      when 1719 => pixel <= "001101";
      when 1720 => pixel <= "001101";
      when 1721 => pixel <= "001101";
      when 1722 => pixel <= "000000";
      when 1723 => pixel <= "000000";
      when 1724 => pixel <= "000000";
      when 1725 => pixel <= "000000";
      when 1726 => pixel <= "000000";
      when 1727 => pixel <= "000000";
      when 1728 => pixel <= "000000";
      when 1729 => pixel <= "000000";
      when 1730 => pixel <= "000000";
      when 1731 => pixel <= "000000";
      when 1732 => pixel <= "000000";
      when 1733 => pixel <= "000000";
      when 1734 => pixel <= "000000";
      when 1735 => pixel <= "000000";
      when 1736 => pixel <= "000000";
      when 1737 => pixel <= "000000";
      when 1738 => pixel <= "000000";
      when 1739 => pixel <= "000000";
      when 1740 => pixel <= "000000";
      when 1741 => pixel <= "000000";
      when 1742 => pixel <= "000000";
      when 1743 => pixel <= "000000";
      when 1744 => pixel <= "000000";
      when 1745 => pixel <= "000000";
      when 1746 => pixel <= "000000";
      when 1747 => pixel <= "000000";
      when 1748 => pixel <= "000000";
      when 1749 => pixel <= "000000";
      when 1750 => pixel <= "000000";
      when 1751 => pixel <= "000000";
      when 1752 => pixel <= "000000";
      when 1753 => pixel <= "000000";
      when 1754 => pixel <= "000000";
      when 1755 => pixel <= "000000";
      when 1756 => pixel <= "000000";
      when 1757 => pixel <= "000000";
      when 1758 => pixel <= "000000";
      when 1759 => pixel <= "000000";
      when 1760 => pixel <= "000000";
      when 1761 => pixel <= "000000";
      when 1762 => pixel <= "000000";
      when 1763 => pixel <= "000000";
      when 1764 => pixel <= "000000";
      when 1765 => pixel <= "000000";
      when 1766 => pixel <= "000000";
      when 1767 => pixel <= "000000";
      when 1768 => pixel <= "000000";
      when 1769 => pixel <= "000000";
      when 1770 => pixel <= "000000";
      when 1771 => pixel <= "000000";
      when 1772 => pixel <= "000000";
      when 1773 => pixel <= "000000";
      when 1774 => pixel <= "000000";
      when 1775 => pixel <= "000000";
      when 1776 => pixel <= "000000";
      when 1777 => pixel <= "000000";
      when 1778 => pixel <= "000000";
      when 1779 => pixel <= "000000";
      when 1780 => pixel <= "000000";
      when 1781 => pixel <= "000000";
      when 1782 => pixel <= "000000";
      when 1783 => pixel <= "000000";
      when 1784 => pixel <= "000000";
      when 1785 => pixel <= "000000";
      when 1786 => pixel <= "000000";
      when 1787 => pixel <= "000000";
      when 1788 => pixel <= "000000";
      when 1789 => pixel <= "000000";
      when 1790 => pixel <= "000000";
      when 1791 => pixel <= "000000";
      when 1792 => pixel <= "000000";
      when 1793 => pixel <= "000000";
      when 1794 => pixel <= "001101";
      when 1795 => pixel <= "001101";
      when 1796 => pixel <= "000000";
      when 1797 => pixel <= "000000";
      when 1798 => pixel <= "000000";
      when 1799 => pixel <= "000000";
      when 1800 => pixel <= "000000";
      when 1801 => pixel <= "000000";
      when 1802 => pixel <= "000000";
      when 1803 => pixel <= "001101";
      when 1804 => pixel <= "001101";
      when 1805 => pixel <= "000000";
      when 1806 => pixel <= "000000";
      when 1807 => pixel <= "000000";
      when 1808 => pixel <= "001101";
      when 1809 => pixel <= "001101";
      when 1810 => pixel <= "000000";
      when 1811 => pixel <= "000000";
      when 1812 => pixel <= "001101";
      when 1813 => pixel <= "001101";
      when 1814 => pixel <= "000000";
      when 1815 => pixel <= "001101";
      when 1816 => pixel <= "000000";
      when 1817 => pixel <= "001101";
      when 1818 => pixel <= "001101";
      when 1819 => pixel <= "000000";
      when 1820 => pixel <= "000000";
      when 1821 => pixel <= "000000";
      when 1822 => pixel <= "001101";
      when 1823 => pixel <= "001101";
      when 1824 => pixel <= "001101";
      when 1825 => pixel <= "001101";
      when 1826 => pixel <= "000000";
      when 1827 => pixel <= "000000";
      when 1828 => pixel <= "000000";
      when 1829 => pixel <= "000000";
      when 1830 => pixel <= "000000";
      when 1831 => pixel <= "000000";
      when 1832 => pixel <= "000000";
      when 1833 => pixel <= "000000";
      when 1834 => pixel <= "000000";
      when 1835 => pixel <= "000000";
      when 1836 => pixel <= "000000";
      when 1837 => pixel <= "000000";
      when 1838 => pixel <= "000000";
      when 1839 => pixel <= "001101";
      when 1840 => pixel <= "001101";
      when 1841 => pixel <= "001101";
      when 1842 => pixel <= "000000";
      when 1843 => pixel <= "000000";
      when 1844 => pixel <= "000000";
      when 1845 => pixel <= "001101";
      when 1846 => pixel <= "001101";
      when 1847 => pixel <= "000000";
      when 1848 => pixel <= "000000";
      when 1849 => pixel <= "001101";
      when 1850 => pixel <= "001101";
      when 1851 => pixel <= "000000";
      when 1852 => pixel <= "000000";
      when 1853 => pixel <= "000000";
      when 1854 => pixel <= "001101";
      when 1855 => pixel <= "001101";
      when 1856 => pixel <= "000000";
      when 1857 => pixel <= "000000";
      when 1858 => pixel <= "000000";
      when 1859 => pixel <= "001101";
      when 1860 => pixel <= "001101";
      when 1861 => pixel <= "001101";
      when 1862 => pixel <= "001101";
      when 1863 => pixel <= "000000";
      when 1864 => pixel <= "000000";
      when 1865 => pixel <= "000000";
      when 1866 => pixel <= "000000";
      when 1867 => pixel <= "000000";
      when 1868 => pixel <= "001101";
      when 1869 => pixel <= "001101";
      when 1870 => pixel <= "001101";
      when 1871 => pixel <= "001101";
      when 1872 => pixel <= "001101";
      when 1873 => pixel <= "000000";
      when 1874 => pixel <= "000000";
      when 1875 => pixel <= "000000";
      when 1876 => pixel <= "000000";
      when 1877 => pixel <= "000000";
      when 1878 => pixel <= "000000";
      when 1879 => pixel <= "001101";
      when 1880 => pixel <= "001101";
      when 1881 => pixel <= "000000";
      when 1882 => pixel <= "000000";
      when 1883 => pixel <= "000000";
      when 1884 => pixel <= "000000";
      when 1885 => pixel <= "000000";
      when 1886 => pixel <= "000000";
      when 1887 => pixel <= "000000";
      when 1888 => pixel <= "000000";
      when 1889 => pixel <= "000000";
      when 1890 => pixel <= "000000";
      when 1891 => pixel <= "000000";
      when 1892 => pixel <= "000000";
      when 1893 => pixel <= "000000";
      when 1894 => pixel <= "000000";
      when 1895 => pixel <= "000000";
      when 1896 => pixel <= "000000";
      when 1897 => pixel <= "000000";
      when 1898 => pixel <= "000000";
      when 1899 => pixel <= "000000";
      when 1900 => pixel <= "000000";
      when 1901 => pixel <= "000000";
      when 1902 => pixel <= "000000";
      when 1903 => pixel <= "000000";
      when 1904 => pixel <= "000000";
      when 1905 => pixel <= "000000";
      when 1906 => pixel <= "000000";
      when 1907 => pixel <= "000000";
      when 1908 => pixel <= "000000";
      when 1909 => pixel <= "000000";
      when 1910 => pixel <= "000000";
      when 1911 => pixel <= "000000";
      when 1912 => pixel <= "000000";
      when 1913 => pixel <= "000000";
      when 1914 => pixel <= "000000";
      when 1915 => pixel <= "000000";
      when 1916 => pixel <= "000000";
      when 1917 => pixel <= "000000";
      when 1918 => pixel <= "000000";
      when 1919 => pixel <= "000000";
      when 1920 => pixel <= "000000";
      when 1921 => pixel <= "000000";
      when 1922 => pixel <= "000000";
      when 1923 => pixel <= "000000";
      when 1924 => pixel <= "000000";
      when 1925 => pixel <= "000000";
      when 1926 => pixel <= "000000";
      when 1927 => pixel <= "000000";
      when 1928 => pixel <= "000000";
      when 1929 => pixel <= "000000";
      when 1930 => pixel <= "000000";
      when 1931 => pixel <= "000000";
      when 1932 => pixel <= "000000";
      when 1933 => pixel <= "000000";
      when 1934 => pixel <= "000000";
      when 1935 => pixel <= "000000";
      when 1936 => pixel <= "000000";
      when 1937 => pixel <= "000000";
      when 1938 => pixel <= "000000";
      when 1939 => pixel <= "000000";
      when 1940 => pixel <= "000000";
      when 1941 => pixel <= "000000";
      when 1942 => pixel <= "000000";
      when 1943 => pixel <= "000000";
      when 1944 => pixel <= "000000";
      when 1945 => pixel <= "000000";
      when 1946 => pixel <= "000000";
      when 1947 => pixel <= "000000";
      when 1948 => pixel <= "000000";
      when 1949 => pixel <= "000000";
      when 1950 => pixel <= "000000";
      when 1951 => pixel <= "000000";
      when 1952 => pixel <= "000000";
      when 1953 => pixel <= "000000";
      when 1954 => pixel <= "001101";
      when 1955 => pixel <= "001101";
      when 1956 => pixel <= "000000";
      when 1957 => pixel <= "001101";
      when 1958 => pixel <= "001101";
      when 1959 => pixel <= "001101";
      when 1960 => pixel <= "001101";
      when 1961 => pixel <= "000000";
      when 1962 => pixel <= "000000";
      when 1963 => pixel <= "001101";
      when 1964 => pixel <= "001101";
      when 1965 => pixel <= "001101";
      when 1966 => pixel <= "001101";
      when 1967 => pixel <= "001101";
      when 1968 => pixel <= "001101";
      when 1969 => pixel <= "001101";
      when 1970 => pixel <= "000000";
      when 1971 => pixel <= "000000";
      when 1972 => pixel <= "001101";
      when 1973 => pixel <= "001101";
      when 1974 => pixel <= "000000";
      when 1975 => pixel <= "000000";
      when 1976 => pixel <= "000000";
      when 1977 => pixel <= "001101";
      when 1978 => pixel <= "001101";
      when 1979 => pixel <= "000000";
      when 1980 => pixel <= "000000";
      when 1981 => pixel <= "000000";
      when 1982 => pixel <= "001101";
      when 1983 => pixel <= "001101";
      when 1984 => pixel <= "000000";
      when 1985 => pixel <= "001101";
      when 1986 => pixel <= "000000";
      when 1987 => pixel <= "000000";
      when 1988 => pixel <= "000000";
      when 1989 => pixel <= "000000";
      when 1990 => pixel <= "000000";
      when 1991 => pixel <= "000000";
      when 1992 => pixel <= "000000";
      when 1993 => pixel <= "000000";
      when 1994 => pixel <= "000000";
      when 1995 => pixel <= "000000";
      when 1996 => pixel <= "000000";
      when 1997 => pixel <= "000000";
      when 1998 => pixel <= "000000";
      when 1999 => pixel <= "001101";
      when 2000 => pixel <= "001101";
      when 2001 => pixel <= "001101";
      when 2002 => pixel <= "000000";
      when 2003 => pixel <= "000000";
      when 2004 => pixel <= "000000";
      when 2005 => pixel <= "001101";
      when 2006 => pixel <= "001101";
      when 2007 => pixel <= "000000";
      when 2008 => pixel <= "000000";
      when 2009 => pixel <= "001101";
      when 2010 => pixel <= "001101";
      when 2011 => pixel <= "000000";
      when 2012 => pixel <= "000000";
      when 2013 => pixel <= "000000";
      when 2014 => pixel <= "001101";
      when 2015 => pixel <= "001101";
      when 2016 => pixel <= "000000";
      when 2017 => pixel <= "000000";
      when 2018 => pixel <= "000000";
      when 2019 => pixel <= "001101";
      when 2020 => pixel <= "001101";
      when 2021 => pixel <= "000000";
      when 2022 => pixel <= "001101";
      when 2023 => pixel <= "000000";
      when 2024 => pixel <= "000000";
      when 2025 => pixel <= "000000";
      when 2026 => pixel <= "000000";
      when 2027 => pixel <= "000000";
      when 2028 => pixel <= "001101";
      when 2029 => pixel <= "001101";
      when 2030 => pixel <= "000000";
      when 2031 => pixel <= "001101";
      when 2032 => pixel <= "001101";
      when 2033 => pixel <= "000000";
      when 2034 => pixel <= "000000";
      when 2035 => pixel <= "000000";
      when 2036 => pixel <= "000000";
      when 2037 => pixel <= "000000";
      when 2038 => pixel <= "000000";
      when 2039 => pixel <= "001101";
      when 2040 => pixel <= "001101";
      when 2041 => pixel <= "000000";
      when 2042 => pixel <= "000000";
      when 2043 => pixel <= "000000";
      when 2044 => pixel <= "000000";
      when 2045 => pixel <= "000000";
      when 2046 => pixel <= "000000";
      when 2047 => pixel <= "000000";
      when 2048 => pixel <= "000000";
      when 2049 => pixel <= "000000";
      when 2050 => pixel <= "000000";
      when 2051 => pixel <= "000000";
      when 2052 => pixel <= "000000";
      when 2053 => pixel <= "000000";
      when 2054 => pixel <= "000000";
      when 2055 => pixel <= "000000";
      when 2056 => pixel <= "000000";
      when 2057 => pixel <= "000000";
      when 2058 => pixel <= "000000";
      when 2059 => pixel <= "000000";
      when 2060 => pixel <= "000000";
      when 2061 => pixel <= "000000";
      when 2062 => pixel <= "000000";
      when 2063 => pixel <= "000000";
      when 2064 => pixel <= "000000";
      when 2065 => pixel <= "000000";
      when 2066 => pixel <= "000000";
      when 2067 => pixel <= "000000";
      when 2068 => pixel <= "000000";
      when 2069 => pixel <= "000000";
      when 2070 => pixel <= "000000";
      when 2071 => pixel <= "000000";
      when 2072 => pixel <= "000000";
      when 2073 => pixel <= "000000";
      when 2074 => pixel <= "000000";
      when 2075 => pixel <= "000000";
      when 2076 => pixel <= "000000";
      when 2077 => pixel <= "000000";
      when 2078 => pixel <= "000000";
      when 2079 => pixel <= "000000";
      when 2080 => pixel <= "000000";
      when 2081 => pixel <= "000000";
      when 2082 => pixel <= "000000";
      when 2083 => pixel <= "000000";
      when 2084 => pixel <= "000000";
      when 2085 => pixel <= "000000";
      when 2086 => pixel <= "000000";
      when 2087 => pixel <= "000000";
      when 2088 => pixel <= "000000";
      when 2089 => pixel <= "000000";
      when 2090 => pixel <= "000000";
      when 2091 => pixel <= "000000";
      when 2092 => pixel <= "000000";
      when 2093 => pixel <= "000000";
      when 2094 => pixel <= "000000";
      when 2095 => pixel <= "000000";
      when 2096 => pixel <= "000000";
      when 2097 => pixel <= "000000";
      when 2098 => pixel <= "000000";
      when 2099 => pixel <= "000000";
      when 2100 => pixel <= "000000";
      when 2101 => pixel <= "000000";
      when 2102 => pixel <= "000000";
      when 2103 => pixel <= "000000";
      when 2104 => pixel <= "000000";
      when 2105 => pixel <= "000000";
      when 2106 => pixel <= "000000";
      when 2107 => pixel <= "000000";
      when 2108 => pixel <= "000000";
      when 2109 => pixel <= "000000";
      when 2110 => pixel <= "000000";
      when 2111 => pixel <= "000000";
      when 2112 => pixel <= "000000";
      when 2113 => pixel <= "000000";
      when 2114 => pixel <= "001101";
      when 2115 => pixel <= "001101";
      when 2116 => pixel <= "000000";
      when 2117 => pixel <= "000000";
      when 2118 => pixel <= "000000";
      when 2119 => pixel <= "001101";
      when 2120 => pixel <= "001101";
      when 2121 => pixel <= "000000";
      when 2122 => pixel <= "000000";
      when 2123 => pixel <= "001101";
      when 2124 => pixel <= "001101";
      when 2125 => pixel <= "000000";
      when 2126 => pixel <= "000000";
      when 2127 => pixel <= "000000";
      when 2128 => pixel <= "001101";
      when 2129 => pixel <= "001101";
      when 2130 => pixel <= "000000";
      when 2131 => pixel <= "000000";
      when 2132 => pixel <= "001101";
      when 2133 => pixel <= "001101";
      when 2134 => pixel <= "000000";
      when 2135 => pixel <= "000000";
      when 2136 => pixel <= "000000";
      when 2137 => pixel <= "001101";
      when 2138 => pixel <= "001101";
      when 2139 => pixel <= "000000";
      when 2140 => pixel <= "000000";
      when 2141 => pixel <= "000000";
      when 2142 => pixel <= "001101";
      when 2143 => pixel <= "001101";
      when 2144 => pixel <= "000000";
      when 2145 => pixel <= "000000";
      when 2146 => pixel <= "000000";
      when 2147 => pixel <= "000000";
      when 2148 => pixel <= "000000";
      when 2149 => pixel <= "000000";
      when 2150 => pixel <= "000000";
      when 2151 => pixel <= "000000";
      when 2152 => pixel <= "000000";
      when 2153 => pixel <= "000000";
      when 2154 => pixel <= "000000";
      when 2155 => pixel <= "000000";
      when 2156 => pixel <= "000000";
      when 2157 => pixel <= "000000";
      when 2158 => pixel <= "000000";
      when 2159 => pixel <= "001101";
      when 2160 => pixel <= "001101";
      when 2161 => pixel <= "001101";
      when 2162 => pixel <= "000000";
      when 2163 => pixel <= "000000";
      when 2164 => pixel <= "000000";
      when 2165 => pixel <= "001101";
      when 2166 => pixel <= "001101";
      when 2167 => pixel <= "000000";
      when 2168 => pixel <= "000000";
      when 2169 => pixel <= "001101";
      when 2170 => pixel <= "001101";
      when 2171 => pixel <= "000000";
      when 2172 => pixel <= "000000";
      when 2173 => pixel <= "000000";
      when 2174 => pixel <= "001101";
      when 2175 => pixel <= "001101";
      when 2176 => pixel <= "000000";
      when 2177 => pixel <= "000000";
      when 2178 => pixel <= "000000";
      when 2179 => pixel <= "001101";
      when 2180 => pixel <= "001101";
      when 2181 => pixel <= "000000";
      when 2182 => pixel <= "000000";
      when 2183 => pixel <= "000000";
      when 2184 => pixel <= "000000";
      when 2185 => pixel <= "000000";
      when 2186 => pixel <= "000000";
      when 2187 => pixel <= "000000";
      when 2188 => pixel <= "001101";
      when 2189 => pixel <= "001101";
      when 2190 => pixel <= "000000";
      when 2191 => pixel <= "000000";
      when 2192 => pixel <= "001101";
      when 2193 => pixel <= "001101";
      when 2194 => pixel <= "000000";
      when 2195 => pixel <= "000000";
      when 2196 => pixel <= "000000";
      when 2197 => pixel <= "000000";
      when 2198 => pixel <= "000000";
      when 2199 => pixel <= "001101";
      when 2200 => pixel <= "001101";
      when 2201 => pixel <= "000000";
      when 2202 => pixel <= "000000";
      when 2203 => pixel <= "000000";
      when 2204 => pixel <= "000000";
      when 2205 => pixel <= "000000";
      when 2206 => pixel <= "000000";
      when 2207 => pixel <= "000000";
      when 2208 => pixel <= "000000";
      when 2209 => pixel <= "000000";
      when 2210 => pixel <= "000000";
      when 2211 => pixel <= "000000";
      when 2212 => pixel <= "000000";
      when 2213 => pixel <= "000000";
      when 2214 => pixel <= "000000";
      when 2215 => pixel <= "000000";
      when 2216 => pixel <= "000000";
      when 2217 => pixel <= "000000";
      when 2218 => pixel <= "000000";
      when 2219 => pixel <= "000000";
      when 2220 => pixel <= "000000";
      when 2221 => pixel <= "000000";
      when 2222 => pixel <= "000000";
      when 2223 => pixel <= "000000";
      when 2224 => pixel <= "000000";
      when 2225 => pixel <= "000000";
      when 2226 => pixel <= "000000";
      when 2227 => pixel <= "000000";
      when 2228 => pixel <= "000000";
      when 2229 => pixel <= "000000";
      when 2230 => pixel <= "000000";
      when 2231 => pixel <= "000000";
      when 2232 => pixel <= "000000";
      when 2233 => pixel <= "000000";
      when 2234 => pixel <= "000000";
      when 2235 => pixel <= "000000";
      when 2236 => pixel <= "000000";
      when 2237 => pixel <= "000000";
      when 2238 => pixel <= "000000";
      when 2239 => pixel <= "000000";
      when 2240 => pixel <= "000000";
      when 2241 => pixel <= "000000";
      when 2242 => pixel <= "000000";
      when 2243 => pixel <= "000000";
      when 2244 => pixel <= "000000";
      when 2245 => pixel <= "000000";
      when 2246 => pixel <= "000000";
      when 2247 => pixel <= "000000";
      when 2248 => pixel <= "000000";
      when 2249 => pixel <= "000000";
      when 2250 => pixel <= "000000";
      when 2251 => pixel <= "000000";
      when 2252 => pixel <= "000000";
      when 2253 => pixel <= "000000";
      when 2254 => pixel <= "000000";
      when 2255 => pixel <= "000000";
      when 2256 => pixel <= "000000";
      when 2257 => pixel <= "000000";
      when 2258 => pixel <= "000000";
      when 2259 => pixel <= "000000";
      when 2260 => pixel <= "000000";
      when 2261 => pixel <= "000000";
      when 2262 => pixel <= "000000";
      when 2263 => pixel <= "000000";
      when 2264 => pixel <= "000000";
      when 2265 => pixel <= "000000";
      when 2266 => pixel <= "000000";
      when 2267 => pixel <= "000000";
      when 2268 => pixel <= "000000";
      when 2269 => pixel <= "000000";
      when 2270 => pixel <= "000000";
      when 2271 => pixel <= "000000";
      when 2272 => pixel <= "000000";
      when 2273 => pixel <= "000000";
      when 2274 => pixel <= "001101";
      when 2275 => pixel <= "001101";
      when 2276 => pixel <= "000000";
      when 2277 => pixel <= "000000";
      when 2278 => pixel <= "000000";
      when 2279 => pixel <= "001101";
      when 2280 => pixel <= "001101";
      when 2281 => pixel <= "000000";
      when 2282 => pixel <= "000000";
      when 2283 => pixel <= "001101";
      when 2284 => pixel <= "001101";
      when 2285 => pixel <= "000000";
      when 2286 => pixel <= "000000";
      when 2287 => pixel <= "000000";
      when 2288 => pixel <= "001101";
      when 2289 => pixel <= "001101";
      when 2290 => pixel <= "000000";
      when 2291 => pixel <= "000000";
      when 2292 => pixel <= "001101";
      when 2293 => pixel <= "001101";
      when 2294 => pixel <= "000000";
      when 2295 => pixel <= "000000";
      when 2296 => pixel <= "000000";
      when 2297 => pixel <= "001101";
      when 2298 => pixel <= "001101";
      when 2299 => pixel <= "000000";
      when 2300 => pixel <= "000000";
      when 2301 => pixel <= "000000";
      when 2302 => pixel <= "001101";
      when 2303 => pixel <= "001101";
      when 2304 => pixel <= "000000";
      when 2305 => pixel <= "000000";
      when 2306 => pixel <= "000000";
      when 2307 => pixel <= "001101";
      when 2308 => pixel <= "000000";
      when 2309 => pixel <= "000000";
      when 2310 => pixel <= "000000";
      when 2311 => pixel <= "000000";
      when 2312 => pixel <= "000000";
      when 2313 => pixel <= "000000";
      when 2314 => pixel <= "000000";
      when 2315 => pixel <= "000000";
      when 2316 => pixel <= "000000";
      when 2317 => pixel <= "000000";
      when 2318 => pixel <= "000000";
      when 2319 => pixel <= "001101";
      when 2320 => pixel <= "001101";
      when 2321 => pixel <= "001101";
      when 2322 => pixel <= "000000";
      when 2323 => pixel <= "000000";
      when 2324 => pixel <= "000000";
      when 2325 => pixel <= "001101";
      when 2326 => pixel <= "001101";
      when 2327 => pixel <= "000000";
      when 2328 => pixel <= "000000";
      when 2329 => pixel <= "000000";
      when 2330 => pixel <= "001101";
      when 2331 => pixel <= "001101";
      when 2332 => pixel <= "000000";
      when 2333 => pixel <= "001101";
      when 2334 => pixel <= "001101";
      when 2335 => pixel <= "000000";
      when 2336 => pixel <= "000000";
      when 2337 => pixel <= "000000";
      when 2338 => pixel <= "000000";
      when 2339 => pixel <= "001101";
      when 2340 => pixel <= "001101";
      when 2341 => pixel <= "000000";
      when 2342 => pixel <= "000000";
      when 2343 => pixel <= "000000";
      when 2344 => pixel <= "001101";
      when 2345 => pixel <= "000000";
      when 2346 => pixel <= "000000";
      when 2347 => pixel <= "000000";
      when 2348 => pixel <= "001101";
      when 2349 => pixel <= "001101";
      when 2350 => pixel <= "000000";
      when 2351 => pixel <= "000000";
      when 2352 => pixel <= "001101";
      when 2353 => pixel <= "001101";
      when 2354 => pixel <= "000000";
      when 2355 => pixel <= "000000";
      when 2356 => pixel <= "000000";
      when 2357 => pixel <= "000000";
      when 2358 => pixel <= "000000";
      when 2359 => pixel <= "000000";
      when 2360 => pixel <= "000000";
      when 2361 => pixel <= "000000";
      when 2362 => pixel <= "000000";
      when 2363 => pixel <= "000000";
      when 2364 => pixel <= "000000";
      when 2365 => pixel <= "000000";
      when 2366 => pixel <= "000000";
      when 2367 => pixel <= "000000";
      when 2368 => pixel <= "000000";
      when 2369 => pixel <= "000000";
      when 2370 => pixel <= "000000";
      when 2371 => pixel <= "000000";
      when 2372 => pixel <= "000000";
      when 2373 => pixel <= "000000";
      when 2374 => pixel <= "000000";
      when 2375 => pixel <= "000000";
      when 2376 => pixel <= "000000";
      when 2377 => pixel <= "000000";
      when 2378 => pixel <= "000000";
      when 2379 => pixel <= "000000";
      when 2380 => pixel <= "000000";
      when 2381 => pixel <= "000000";
      when 2382 => pixel <= "000000";
      when 2383 => pixel <= "000000";
      when 2384 => pixel <= "000000";
      when 2385 => pixel <= "000000";
      when 2386 => pixel <= "000000";
      when 2387 => pixel <= "000000";
      when 2388 => pixel <= "000000";
      when 2389 => pixel <= "000000";
      when 2390 => pixel <= "000000";
      when 2391 => pixel <= "000000";
      when 2392 => pixel <= "000000";
      when 2393 => pixel <= "000000";
      when 2394 => pixel <= "000000";
      when 2395 => pixel <= "000000";
      when 2396 => pixel <= "000000";
      when 2397 => pixel <= "000000";
      when 2398 => pixel <= "000000";
      when 2399 => pixel <= "000000";
      when 2400 => pixel <= "000000";
      when 2401 => pixel <= "000000";
      when 2402 => pixel <= "000000";
      when 2403 => pixel <= "000000";
      when 2404 => pixel <= "000000";
      when 2405 => pixel <= "000000";
      when 2406 => pixel <= "000000";
      when 2407 => pixel <= "000000";
      when 2408 => pixel <= "000000";
      when 2409 => pixel <= "000000";
      when 2410 => pixel <= "000000";
      when 2411 => pixel <= "000000";
      when 2412 => pixel <= "000000";
      when 2413 => pixel <= "000000";
      when 2414 => pixel <= "000000";
      when 2415 => pixel <= "000000";
      when 2416 => pixel <= "000000";
      when 2417 => pixel <= "000000";
      when 2418 => pixel <= "000000";
      when 2419 => pixel <= "000000";
      when 2420 => pixel <= "000000";
      when 2421 => pixel <= "000000";
      when 2422 => pixel <= "000000";
      when 2423 => pixel <= "000000";
      when 2424 => pixel <= "000000";
      when 2425 => pixel <= "000000";
      when 2426 => pixel <= "000000";
      when 2427 => pixel <= "000000";
      when 2428 => pixel <= "000000";
      when 2429 => pixel <= "000000";
      when 2430 => pixel <= "000000";
      when 2431 => pixel <= "000000";
      when 2432 => pixel <= "000000";
      when 2433 => pixel <= "000000";
      when 2434 => pixel <= "000000";
      when 2435 => pixel <= "001101";
      when 2436 => pixel <= "001101";
      when 2437 => pixel <= "000000";
      when 2438 => pixel <= "000000";
      when 2439 => pixel <= "001101";
      when 2440 => pixel <= "001101";
      when 2441 => pixel <= "000000";
      when 2442 => pixel <= "000000";
      when 2443 => pixel <= "001101";
      when 2444 => pixel <= "001101";
      when 2445 => pixel <= "000000";
      when 2446 => pixel <= "000000";
      when 2447 => pixel <= "000000";
      when 2448 => pixel <= "001101";
      when 2449 => pixel <= "001101";
      when 2450 => pixel <= "000000";
      when 2451 => pixel <= "000000";
      when 2452 => pixel <= "001101";
      when 2453 => pixel <= "001101";
      when 2454 => pixel <= "000000";
      when 2455 => pixel <= "000000";
      when 2456 => pixel <= "000000";
      when 2457 => pixel <= "001101";
      when 2458 => pixel <= "001101";
      when 2459 => pixel <= "000000";
      when 2460 => pixel <= "000000";
      when 2461 => pixel <= "000000";
      when 2462 => pixel <= "001101";
      when 2463 => pixel <= "001101";
      when 2464 => pixel <= "000000";
      when 2465 => pixel <= "000000";
      when 2466 => pixel <= "001101";
      when 2467 => pixel <= "001101";
      when 2468 => pixel <= "000000";
      when 2469 => pixel <= "000000";
      when 2470 => pixel <= "000000";
      when 2471 => pixel <= "000000";
      when 2472 => pixel <= "000000";
      when 2473 => pixel <= "000000";
      when 2474 => pixel <= "000000";
      when 2475 => pixel <= "000000";
      when 2476 => pixel <= "000000";
      when 2477 => pixel <= "000000";
      when 2478 => pixel <= "000000";
      when 2479 => pixel <= "001101";
      when 2480 => pixel <= "001101";
      when 2481 => pixel <= "001101";
      when 2482 => pixel <= "000000";
      when 2483 => pixel <= "000000";
      when 2484 => pixel <= "000000";
      when 2485 => pixel <= "001101";
      when 2486 => pixel <= "001101";
      when 2487 => pixel <= "000000";
      when 2488 => pixel <= "000000";
      when 2489 => pixel <= "000000";
      when 2490 => pixel <= "000000";
      when 2491 => pixel <= "001101";
      when 2492 => pixel <= "001101";
      when 2493 => pixel <= "001101";
      when 2494 => pixel <= "000000";
      when 2495 => pixel <= "000000";
      when 2496 => pixel <= "000000";
      when 2497 => pixel <= "000000";
      when 2498 => pixel <= "000000";
      when 2499 => pixel <= "001101";
      when 2500 => pixel <= "001101";
      when 2501 => pixel <= "000000";
      when 2502 => pixel <= "000000";
      when 2503 => pixel <= "001101";
      when 2504 => pixel <= "001101";
      when 2505 => pixel <= "000000";
      when 2506 => pixel <= "000000";
      when 2507 => pixel <= "000000";
      when 2508 => pixel <= "001101";
      when 2509 => pixel <= "001101";
      when 2510 => pixel <= "000000";
      when 2511 => pixel <= "000000";
      when 2512 => pixel <= "001101";
      when 2513 => pixel <= "001101";
      when 2514 => pixel <= "000000";
      when 2515 => pixel <= "000000";
      when 2516 => pixel <= "000000";
      when 2517 => pixel <= "000000";
      when 2518 => pixel <= "000000";
      when 2519 => pixel <= "001101";
      when 2520 => pixel <= "001101";
      when 2521 => pixel <= "000000";
      when 2522 => pixel <= "000000";
      when 2523 => pixel <= "000000";
      when 2524 => pixel <= "000000";
      when 2525 => pixel <= "000000";
      when 2526 => pixel <= "000000";
      when 2527 => pixel <= "000000";
      when 2528 => pixel <= "000000";
      when 2529 => pixel <= "000000";
      when 2530 => pixel <= "000000";
      when 2531 => pixel <= "000000";
      when 2532 => pixel <= "000000";
      when 2533 => pixel <= "000000";
      when 2534 => pixel <= "000000";
      when 2535 => pixel <= "000000";
      when 2536 => pixel <= "000000";
      when 2537 => pixel <= "000000";
      when 2538 => pixel <= "000000";
      when 2539 => pixel <= "000000";
      when 2540 => pixel <= "000000";
      when 2541 => pixel <= "000000";
      when 2542 => pixel <= "000000";
      when 2543 => pixel <= "000000";
      when 2544 => pixel <= "000000";
      when 2545 => pixel <= "000000";
      when 2546 => pixel <= "000000";
      when 2547 => pixel <= "000000";
      when 2548 => pixel <= "000000";
      when 2549 => pixel <= "000000";
      when 2550 => pixel <= "000000";
      when 2551 => pixel <= "000000";
      when 2552 => pixel <= "000000";
      when 2553 => pixel <= "000000";
      when 2554 => pixel <= "000000";
      when 2555 => pixel <= "000000";
      when 2556 => pixel <= "000000";
      when 2557 => pixel <= "000000";
      when 2558 => pixel <= "000000";
      when 2559 => pixel <= "000000";
      when 2560 => pixel <= "000000";
      when 2561 => pixel <= "000000";
      when 2562 => pixel <= "000000";
      when 2563 => pixel <= "000000";
      when 2564 => pixel <= "000000";
      when 2565 => pixel <= "000000";
      when 2566 => pixel <= "000000";
      when 2567 => pixel <= "000000";
      when 2568 => pixel <= "000000";
      when 2569 => pixel <= "000000";
      when 2570 => pixel <= "000000";
      when 2571 => pixel <= "000000";
      when 2572 => pixel <= "000000";
      when 2573 => pixel <= "000000";
      when 2574 => pixel <= "000000";
      when 2575 => pixel <= "000000";
      when 2576 => pixel <= "000000";
      when 2577 => pixel <= "000000";
      when 2578 => pixel <= "000000";
      when 2579 => pixel <= "000000";
      when 2580 => pixel <= "000000";
      when 2581 => pixel <= "000000";
      when 2582 => pixel <= "000000";
      when 2583 => pixel <= "000000";
      when 2584 => pixel <= "000000";
      when 2585 => pixel <= "000000";
      when 2586 => pixel <= "000000";
      when 2587 => pixel <= "000000";
      when 2588 => pixel <= "000000";
      when 2589 => pixel <= "000000";
      when 2590 => pixel <= "000000";
      when 2591 => pixel <= "000000";
      when 2592 => pixel <= "000000";
      when 2593 => pixel <= "000000";
      when 2594 => pixel <= "000000";
      when 2595 => pixel <= "000000";
      when 2596 => pixel <= "001101";
      when 2597 => pixel <= "001101";
      when 2598 => pixel <= "001101";
      when 2599 => pixel <= "000000";
      when 2600 => pixel <= "001101";
      when 2601 => pixel <= "000000";
      when 2602 => pixel <= "000000";
      when 2603 => pixel <= "001101";
      when 2604 => pixel <= "001101";
      when 2605 => pixel <= "000000";
      when 2606 => pixel <= "000000";
      when 2607 => pixel <= "000000";
      when 2608 => pixel <= "001101";
      when 2609 => pixel <= "001101";
      when 2610 => pixel <= "000000";
      when 2611 => pixel <= "000000";
      when 2612 => pixel <= "001101";
      when 2613 => pixel <= "001101";
      when 2614 => pixel <= "000000";
      when 2615 => pixel <= "000000";
      when 2616 => pixel <= "000000";
      when 2617 => pixel <= "001101";
      when 2618 => pixel <= "001101";
      when 2619 => pixel <= "000000";
      when 2620 => pixel <= "000000";
      when 2621 => pixel <= "001101";
      when 2622 => pixel <= "001101";
      when 2623 => pixel <= "001101";
      when 2624 => pixel <= "001101";
      when 2625 => pixel <= "001101";
      when 2626 => pixel <= "001101";
      when 2627 => pixel <= "001101";
      when 2628 => pixel <= "000000";
      when 2629 => pixel <= "000000";
      when 2630 => pixel <= "000000";
      when 2631 => pixel <= "000000";
      when 2632 => pixel <= "000000";
      when 2633 => pixel <= "000000";
      when 2634 => pixel <= "000000";
      when 2635 => pixel <= "000000";
      when 2636 => pixel <= "000000";
      when 2637 => pixel <= "000000";
      when 2638 => pixel <= "000000";
      when 2639 => pixel <= "000000";
      when 2640 => pixel <= "000000";
      when 2641 => pixel <= "001101";
      when 2642 => pixel <= "001101";
      when 2643 => pixel <= "001101";
      when 2644 => pixel <= "001101";
      when 2645 => pixel <= "001101";
      when 2646 => pixel <= "000000";
      when 2647 => pixel <= "000000";
      when 2648 => pixel <= "000000";
      when 2649 => pixel <= "000000";
      when 2650 => pixel <= "000000";
      when 2651 => pixel <= "000000";
      when 2652 => pixel <= "001101";
      when 2653 => pixel <= "000000";
      when 2654 => pixel <= "000000";
      when 2655 => pixel <= "000000";
      when 2656 => pixel <= "000000";
      when 2657 => pixel <= "000000";
      when 2658 => pixel <= "001101";
      when 2659 => pixel <= "001101";
      when 2660 => pixel <= "001101";
      when 2661 => pixel <= "001101";
      when 2662 => pixel <= "001101";
      when 2663 => pixel <= "001101";
      when 2664 => pixel <= "001101";
      when 2665 => pixel <= "000000";
      when 2666 => pixel <= "000000";
      when 2667 => pixel <= "001101";
      when 2668 => pixel <= "001101";
      when 2669 => pixel <= "001101";
      when 2670 => pixel <= "000000";
      when 2671 => pixel <= "000000";
      when 2672 => pixel <= "001101";
      when 2673 => pixel <= "001101";
      when 2674 => pixel <= "000000";
      when 2675 => pixel <= "000000";
      when 2676 => pixel <= "000000";
      when 2677 => pixel <= "000000";
      when 2678 => pixel <= "000000";
      when 2679 => pixel <= "001101";
      when 2680 => pixel <= "001101";
      when 2681 => pixel <= "000000";
      when 2682 => pixel <= "000000";
      when 2683 => pixel <= "000000";
      when 2684 => pixel <= "000000";
      when 2685 => pixel <= "000000";
      when 2686 => pixel <= "000000";
      when 2687 => pixel <= "000000";
      when 2688 => pixel <= "000000";
      when 2689 => pixel <= "000000";
      when 2690 => pixel <= "000000";
      when 2691 => pixel <= "000000";
      when 2692 => pixel <= "000000";
      when 2693 => pixel <= "000000";
      when 2694 => pixel <= "000000";
      when 2695 => pixel <= "000000";
      when 2696 => pixel <= "000000";
      when 2697 => pixel <= "000000";
      when 2698 => pixel <= "000000";
      when 2699 => pixel <= "000000";
      when 2700 => pixel <= "000000";
      when 2701 => pixel <= "000000";
      when 2702 => pixel <= "000000";
      when 2703 => pixel <= "000000";
      when 2704 => pixel <= "000000";
      when 2705 => pixel <= "000000";
      when 2706 => pixel <= "000000";
      when 2707 => pixel <= "000000";
      when 2708 => pixel <= "000000";
      when 2709 => pixel <= "000000";
      when 2710 => pixel <= "000000";
      when 2711 => pixel <= "000000";
      when 2712 => pixel <= "000000";
      when 2713 => pixel <= "000000";
      when 2714 => pixel <= "000000";
      when 2715 => pixel <= "000000";
      when 2716 => pixel <= "000000";
      when 2717 => pixel <= "000000";
      when 2718 => pixel <= "000000";
      when 2719 => pixel <= "000000";
      when 2720 => pixel <= "000000";
      when 2721 => pixel <= "000000";
      when 2722 => pixel <= "000000";
      when 2723 => pixel <= "000000";
      when 2724 => pixel <= "000000";
      when 2725 => pixel <= "000000";
      when 2726 => pixel <= "000000";
      when 2727 => pixel <= "000000";
      when 2728 => pixel <= "000000";
      when 2729 => pixel <= "000000";
      when 2730 => pixel <= "000000";
      when 2731 => pixel <= "000000";
      when 2732 => pixel <= "000000";
      when 2733 => pixel <= "000000";
      when 2734 => pixel <= "000000";
      when 2735 => pixel <= "000000";
      when 2736 => pixel <= "000000";
      when 2737 => pixel <= "000000";
      when 2738 => pixel <= "000000";
      when 2739 => pixel <= "000000";
      when 2740 => pixel <= "000000";
      when 2741 => pixel <= "000000";
      when 2742 => pixel <= "000000";
      when 2743 => pixel <= "000000";
      when 2744 => pixel <= "000000";
      when 2745 => pixel <= "000000";
      when 2746 => pixel <= "000000";
      when 2747 => pixel <= "000000";
      when 2748 => pixel <= "000000";
      when 2749 => pixel <= "000000";
      when 2750 => pixel <= "000000";
      when 2751 => pixel <= "000000";
      when 2752 => pixel <= "000000";
      when 2753 => pixel <= "000000";
      when 2754 => pixel <= "000000";
      when 2755 => pixel <= "000000";
      when 2756 => pixel <= "000000";
      when 2757 => pixel <= "000000";
      when 2758 => pixel <= "000000";
      when 2759 => pixel <= "000000";
      when 2760 => pixel <= "000000";
      when 2761 => pixel <= "000000";
      when 2762 => pixel <= "000000";
      when 2763 => pixel <= "000000";
      when 2764 => pixel <= "000000";
      when 2765 => pixel <= "000000";
      when 2766 => pixel <= "000000";
      when 2767 => pixel <= "000000";
      when 2768 => pixel <= "000000";
      when 2769 => pixel <= "000000";
      when 2770 => pixel <= "000000";
      when 2771 => pixel <= "000000";
      when 2772 => pixel <= "000000";
      when 2773 => pixel <= "000000";
      when 2774 => pixel <= "000000";
      when 2775 => pixel <= "000000";
      when 2776 => pixel <= "000000";
      when 2777 => pixel <= "000000";
      when 2778 => pixel <= "000000";
      when 2779 => pixel <= "000000";
      when 2780 => pixel <= "000000";
      when 2781 => pixel <= "000000";
      when 2782 => pixel <= "000000";
      when 2783 => pixel <= "000000";
      when 2784 => pixel <= "000000";
      when 2785 => pixel <= "000000";
      when 2786 => pixel <= "000000";
      when 2787 => pixel <= "000000";
      when 2788 => pixel <= "000000";
      when 2789 => pixel <= "000000";
      when 2790 => pixel <= "000000";
      when 2791 => pixel <= "000000";
      when 2792 => pixel <= "000000";
      when 2793 => pixel <= "000000";
      when 2794 => pixel <= "000000";
      when 2795 => pixel <= "000000";
      when 2796 => pixel <= "000000";
      when 2797 => pixel <= "000000";
      when 2798 => pixel <= "000000";
      when 2799 => pixel <= "000000";
      when 2800 => pixel <= "000000";
      when 2801 => pixel <= "000000";
      when 2802 => pixel <= "000000";
      when 2803 => pixel <= "000000";
      when 2804 => pixel <= "000000";
      when 2805 => pixel <= "000000";
      when 2806 => pixel <= "000000";
      when 2807 => pixel <= "000000";
      when 2808 => pixel <= "000000";
      when 2809 => pixel <= "000000";
      when 2810 => pixel <= "000000";
      when 2811 => pixel <= "000000";
      when 2812 => pixel <= "000000";
      when 2813 => pixel <= "000000";
      when 2814 => pixel <= "000000";
      when 2815 => pixel <= "000000";
      when 2816 => pixel <= "000000";
      when 2817 => pixel <= "000000";
      when 2818 => pixel <= "000000";
      when 2819 => pixel <= "000000";
      when 2820 => pixel <= "000000";
      when 2821 => pixel <= "000000";
      when 2822 => pixel <= "000000";
      when 2823 => pixel <= "000000";
      when 2824 => pixel <= "000000";
      when 2825 => pixel <= "000000";
      when 2826 => pixel <= "000000";
      when 2827 => pixel <= "000000";
      when 2828 => pixel <= "000000";
      when 2829 => pixel <= "000000";
      when 2830 => pixel <= "000000";
      when 2831 => pixel <= "000000";
      when 2832 => pixel <= "000000";
      when 2833 => pixel <= "000000";
      when 2834 => pixel <= "000000";
      when 2835 => pixel <= "000000";
      when 2836 => pixel <= "000000";
      when 2837 => pixel <= "000000";
      when 2838 => pixel <= "000000";
      when 2839 => pixel <= "000000";
      when 2840 => pixel <= "000000";
      when 2841 => pixel <= "000000";
      when 2842 => pixel <= "000000";
      when 2843 => pixel <= "000000";
      when 2844 => pixel <= "000000";
      when 2845 => pixel <= "000000";
      when 2846 => pixel <= "000000";
      when 2847 => pixel <= "000000";
      when 2848 => pixel <= "000000";
      when 2849 => pixel <= "000000";
      when 2850 => pixel <= "000000";
      when 2851 => pixel <= "000000";
      when 2852 => pixel <= "000000";
      when 2853 => pixel <= "000000";
      when 2854 => pixel <= "000000";
      when 2855 => pixel <= "000000";
      when 2856 => pixel <= "000000";
      when 2857 => pixel <= "000000";
      when 2858 => pixel <= "000000";
      when 2859 => pixel <= "000000";
      when 2860 => pixel <= "000000";
      when 2861 => pixel <= "000000";
      when 2862 => pixel <= "000000";
      when 2863 => pixel <= "000000";
      when 2864 => pixel <= "000000";
      when 2865 => pixel <= "000000";
      when 2866 => pixel <= "000000";
      when 2867 => pixel <= "000000";
      when 2868 => pixel <= "000000";
      when 2869 => pixel <= "000000";
      when 2870 => pixel <= "000000";
      when 2871 => pixel <= "000000";
      when 2872 => pixel <= "000000";
      when 2873 => pixel <= "000000";
      when 2874 => pixel <= "000000";
      when 2875 => pixel <= "000000";
      when 2876 => pixel <= "000000";
      when 2877 => pixel <= "000000";
      when 2878 => pixel <= "000000";
      when 2879 => pixel <= "000000";
      when 2880 => pixel <= "000000";
      when 2881 => pixel <= "000000";
      when 2882 => pixel <= "000000";
      when 2883 => pixel <= "000000";
      when 2884 => pixel <= "000000";
      when 2885 => pixel <= "000000";
      when 2886 => pixel <= "000000";
      when 2887 => pixel <= "000000";
      when 2888 => pixel <= "000000";
      when 2889 => pixel <= "000000";
      when 2890 => pixel <= "000000";
      when 2891 => pixel <= "000000";
      when 2892 => pixel <= "000000";
      when 2893 => pixel <= "000000";
      when 2894 => pixel <= "000000";
      when 2895 => pixel <= "000000";
      when 2896 => pixel <= "000000";
      when 2897 => pixel <= "000000";
      when 2898 => pixel <= "000000";
      when 2899 => pixel <= "000000";
      when 2900 => pixel <= "000000";
      when 2901 => pixel <= "000000";
      when 2902 => pixel <= "000000";
      when 2903 => pixel <= "000000";
      when 2904 => pixel <= "000000";
      when 2905 => pixel <= "000000";
      when 2906 => pixel <= "000000";
      when 2907 => pixel <= "000000";
      when 2908 => pixel <= "000000";
      when 2909 => pixel <= "000000";
      when 2910 => pixel <= "000000";
      when 2911 => pixel <= "000000";
      when 2912 => pixel <= "000000";
      when 2913 => pixel <= "000000";
      when 2914 => pixel <= "000000";
      when 2915 => pixel <= "000000";
      when 2916 => pixel <= "000000";
      when 2917 => pixel <= "000000";
      when 2918 => pixel <= "000000";
      when 2919 => pixel <= "000000";
      when 2920 => pixel <= "000000";
      when 2921 => pixel <= "000000";
      when 2922 => pixel <= "000000";
      when 2923 => pixel <= "000000";
      when 2924 => pixel <= "000000";
      when 2925 => pixel <= "000000";
      when 2926 => pixel <= "000000";
      when 2927 => pixel <= "000000";
      when 2928 => pixel <= "000000";
      when 2929 => pixel <= "000000";
      when 2930 => pixel <= "000000";
      when 2931 => pixel <= "000000";
      when 2932 => pixel <= "000000";
      when 2933 => pixel <= "000000";
      when 2934 => pixel <= "000000";
      when 2935 => pixel <= "000000";
      when 2936 => pixel <= "000000";
      when 2937 => pixel <= "000000";
      when 2938 => pixel <= "000000";
      when 2939 => pixel <= "000000";
      when 2940 => pixel <= "000000";
      when 2941 => pixel <= "000000";
      when 2942 => pixel <= "000000";
      when 2943 => pixel <= "000000";
      when 2944 => pixel <= "000000";
      when 2945 => pixel <= "000000";
      when 2946 => pixel <= "000000";
      when 2947 => pixel <= "000000";
      when 2948 => pixel <= "000000";
      when 2949 => pixel <= "000000";
      when 2950 => pixel <= "000000";
      when 2951 => pixel <= "000000";
      when 2952 => pixel <= "000000";
      when 2953 => pixel <= "000000";
      when 2954 => pixel <= "000000";
      when 2955 => pixel <= "000000";
      when 2956 => pixel <= "000000";
      when 2957 => pixel <= "000000";
      when 2958 => pixel <= "000000";
      when 2959 => pixel <= "000000";
      when 2960 => pixel <= "000000";
      when 2961 => pixel <= "000000";
      when 2962 => pixel <= "000000";
      when 2963 => pixel <= "000000";
      when 2964 => pixel <= "000000";
      when 2965 => pixel <= "000000";
      when 2966 => pixel <= "000000";
      when 2967 => pixel <= "000000";
      when 2968 => pixel <= "000000";
      when 2969 => pixel <= "000000";
      when 2970 => pixel <= "000000";
      when 2971 => pixel <= "000000";
      when 2972 => pixel <= "000000";
      when 2973 => pixel <= "000000";
      when 2974 => pixel <= "000000";
      when 2975 => pixel <= "000000";
      when 2976 => pixel <= "000000";
      when 2977 => pixel <= "000000";
      when 2978 => pixel <= "000000";
      when 2979 => pixel <= "000000";
      when 2980 => pixel <= "000000";
      when 2981 => pixel <= "000000";
      when 2982 => pixel <= "000000";
      when 2983 => pixel <= "000000";
      when 2984 => pixel <= "000000";
      when 2985 => pixel <= "000000";
      when 2986 => pixel <= "000000";
      when 2987 => pixel <= "000000";
      when 2988 => pixel <= "000000";
      when 2989 => pixel <= "000000";
      when 2990 => pixel <= "000000";
      when 2991 => pixel <= "000000";
      when 2992 => pixel <= "000000";
      when 2993 => pixel <= "000000";
      when 2994 => pixel <= "000000";
      when 2995 => pixel <= "000000";
      when 2996 => pixel <= "000000";
      when 2997 => pixel <= "000000";
      when 2998 => pixel <= "000000";
      when 2999 => pixel <= "000000";
      when 3000 => pixel <= "000000";
      when 3001 => pixel <= "000000";
      when 3002 => pixel <= "000000";
      when 3003 => pixel <= "000000";
      when 3004 => pixel <= "000000";
      when 3005 => pixel <= "000000";
      when 3006 => pixel <= "000000";
      when 3007 => pixel <= "000000";
      when 3008 => pixel <= "000000";
      when 3009 => pixel <= "000000";
      when 3010 => pixel <= "000000";
      when 3011 => pixel <= "000000";
      when 3012 => pixel <= "000000";
      when 3013 => pixel <= "000000";
      when 3014 => pixel <= "000000";
      when 3015 => pixel <= "000000";
      when 3016 => pixel <= "000000";
      when 3017 => pixel <= "000000";
      when 3018 => pixel <= "000000";
      when 3019 => pixel <= "000000";
      when 3020 => pixel <= "000000";
      when 3021 => pixel <= "000000";
      when 3022 => pixel <= "000000";
      when 3023 => pixel <= "000000";
      when 3024 => pixel <= "000000";
      when 3025 => pixel <= "000000";
      when 3026 => pixel <= "000000";
      when 3027 => pixel <= "000000";
      when 3028 => pixel <= "000000";
      when 3029 => pixel <= "000000";
      when 3030 => pixel <= "000000";
      when 3031 => pixel <= "000000";
      when 3032 => pixel <= "000000";
      when 3033 => pixel <= "000000";
      when 3034 => pixel <= "000000";
      when 3035 => pixel <= "000000";
      when 3036 => pixel <= "000000";
      when 3037 => pixel <= "000000";
      when 3038 => pixel <= "000000";
      when 3039 => pixel <= "000000";
      when 3040 => pixel <= "000000";
      when 3041 => pixel <= "000000";
      when 3042 => pixel <= "000000";
      when 3043 => pixel <= "000000";
      when 3044 => pixel <= "000000";
      when 3045 => pixel <= "000000";
      when 3046 => pixel <= "000000";
      when 3047 => pixel <= "000000";
      when 3048 => pixel <= "000000";
      when 3049 => pixel <= "000000";
      when 3050 => pixel <= "000000";
      when 3051 => pixel <= "000000";
      when 3052 => pixel <= "000000";
      when 3053 => pixel <= "000000";
      when 3054 => pixel <= "000000";
      when 3055 => pixel <= "000000";
      when 3056 => pixel <= "000000";
      when 3057 => pixel <= "000000";
      when 3058 => pixel <= "000000";
      when 3059 => pixel <= "000000";
      when 3060 => pixel <= "000000";
      when 3061 => pixel <= "000000";
      when 3062 => pixel <= "000000";
      when 3063 => pixel <= "000000";
      when 3064 => pixel <= "000000";
      when 3065 => pixel <= "000000";
      when 3066 => pixel <= "000000";
      when 3067 => pixel <= "000000";
      when 3068 => pixel <= "000000";
      when 3069 => pixel <= "000000";
      when 3070 => pixel <= "000000";
      when 3071 => pixel <= "000000";
      when 3072 => pixel <= "000000";
      when 3073 => pixel <= "000000";
      when 3074 => pixel <= "000000";
      when 3075 => pixel <= "000000";
      when 3076 => pixel <= "000000";
      when 3077 => pixel <= "000000";
      when 3078 => pixel <= "000000";
      when 3079 => pixel <= "000000";
      when 3080 => pixel <= "000000";
      when 3081 => pixel <= "000000";
      when 3082 => pixel <= "000000";
      when 3083 => pixel <= "000000";
      when 3084 => pixel <= "000000";
      when 3085 => pixel <= "000000";
      when 3086 => pixel <= "000000";
      when 3087 => pixel <= "000000";
      when 3088 => pixel <= "000000";
      when 3089 => pixel <= "000000";
      when 3090 => pixel <= "000000";
      when 3091 => pixel <= "000000";
      when 3092 => pixel <= "000000";
      when 3093 => pixel <= "000000";
      when 3094 => pixel <= "000000";
      when 3095 => pixel <= "000000";
      when 3096 => pixel <= "000000";
      when 3097 => pixel <= "000000";
      when 3098 => pixel <= "000000";
      when 3099 => pixel <= "000000";
      when 3100 => pixel <= "000000";
      when 3101 => pixel <= "000000";
      when 3102 => pixel <= "000000";
      when 3103 => pixel <= "000000";
      when 3104 => pixel <= "000000";
      when 3105 => pixel <= "000000";
      when 3106 => pixel <= "000000";
      when 3107 => pixel <= "000000";
      when 3108 => pixel <= "000000";
      when 3109 => pixel <= "000000";
      when 3110 => pixel <= "000000";
      when 3111 => pixel <= "000000";
      when 3112 => pixel <= "000000";
      when 3113 => pixel <= "000000";
      when 3114 => pixel <= "000000";
      when 3115 => pixel <= "000000";
      when 3116 => pixel <= "000000";
      when 3117 => pixel <= "000000";
      when 3118 => pixel <= "000000";
      when 3119 => pixel <= "000000";
      when 3120 => pixel <= "000000";
      when 3121 => pixel <= "000000";
      when 3122 => pixel <= "000000";
      when 3123 => pixel <= "000000";
      when 3124 => pixel <= "000000";
      when 3125 => pixel <= "000000";
      when 3126 => pixel <= "000000";
      when 3127 => pixel <= "000000";
      when 3128 => pixel <= "000000";
      when 3129 => pixel <= "000000";
      when 3130 => pixel <= "000000";
      when 3131 => pixel <= "000000";
      when 3132 => pixel <= "000000";
      when 3133 => pixel <= "000000";
      when 3134 => pixel <= "000000";
      when 3135 => pixel <= "000000";
      when 3136 => pixel <= "000000";
      when 3137 => pixel <= "000000";
      when 3138 => pixel <= "000000";
      when 3139 => pixel <= "000000";
      when 3140 => pixel <= "000000";
      when 3141 => pixel <= "000000";
      when 3142 => pixel <= "000000";
      when 3143 => pixel <= "000000";
      when 3144 => pixel <= "000000";
      when 3145 => pixel <= "000000";
      when 3146 => pixel <= "000000";
      when 3147 => pixel <= "000000";
      when 3148 => pixel <= "000000";
      when 3149 => pixel <= "000000";
      when 3150 => pixel <= "000000";
      when 3151 => pixel <= "000000";
      when 3152 => pixel <= "000000";
      when 3153 => pixel <= "000000";
      when 3154 => pixel <= "000000";
      when 3155 => pixel <= "000000";
      when 3156 => pixel <= "000000";
      when 3157 => pixel <= "000000";
      when 3158 => pixel <= "000000";
      when 3159 => pixel <= "000000";
      when 3160 => pixel <= "000000";
      when 3161 => pixel <= "000000";
      when 3162 => pixel <= "000000";
      when 3163 => pixel <= "000000";
      when 3164 => pixel <= "000000";
      when 3165 => pixel <= "000000";
      when 3166 => pixel <= "000000";
      when 3167 => pixel <= "000000";
      when 3168 => pixel <= "000000";
      when 3169 => pixel <= "000000";
      when 3170 => pixel <= "000000";
      when 3171 => pixel <= "000000";
      when 3172 => pixel <= "000000";
      when 3173 => pixel <= "000000";
      when 3174 => pixel <= "000000";
      when 3175 => pixel <= "000000";
      when 3176 => pixel <= "000000";
      when 3177 => pixel <= "000000";
      when 3178 => pixel <= "000000";
      when 3179 => pixel <= "000000";
      when 3180 => pixel <= "000000";
      when 3181 => pixel <= "000000";
      when 3182 => pixel <= "000000";
      when 3183 => pixel <= "000000";
      when 3184 => pixel <= "000000";
      when 3185 => pixel <= "000000";
      when 3186 => pixel <= "000000";
      when 3187 => pixel <= "000000";
      when 3188 => pixel <= "000000";
      when 3189 => pixel <= "000000";
      when 3190 => pixel <= "000000";
      when 3191 => pixel <= "000000";
      when 3192 => pixel <= "000000";
      when 3193 => pixel <= "000000";
      when 3194 => pixel <= "000000";
      when 3195 => pixel <= "000000";
      when 3196 => pixel <= "000000";
      when 3197 => pixel <= "000000";
      when 3198 => pixel <= "000000";
      when 3199 => pixel <= "000000";
      when 3200 => pixel <= "000000";
      when 3201 => pixel <= "000000";
      when 3202 => pixel <= "000000";
      when 3203 => pixel <= "000000";
      when 3204 => pixel <= "000000";
      when 3205 => pixel <= "000000";
      when 3206 => pixel <= "000000";
      when 3207 => pixel <= "000000";
      when 3208 => pixel <= "000000";
      when 3209 => pixel <= "000000";
      when 3210 => pixel <= "000000";
      when 3211 => pixel <= "000000";
      when 3212 => pixel <= "000000";
      when 3213 => pixel <= "000000";
      when 3214 => pixel <= "000000";
      when 3215 => pixel <= "000000";
      when 3216 => pixel <= "000000";
      when 3217 => pixel <= "000000";
      when 3218 => pixel <= "000000";
      when 3219 => pixel <= "000000";
      when 3220 => pixel <= "000000";
      when 3221 => pixel <= "000000";
      when 3222 => pixel <= "000000";
      when 3223 => pixel <= "000000";
      when 3224 => pixel <= "000000";
      when 3225 => pixel <= "000000";
      when 3226 => pixel <= "000000";
      when 3227 => pixel <= "000000";
      when 3228 => pixel <= "000000";
      when 3229 => pixel <= "000000";
      when 3230 => pixel <= "000000";
      when 3231 => pixel <= "000000";
      when 3232 => pixel <= "000000";
      when 3233 => pixel <= "000000";
      when 3234 => pixel <= "000000";
      when 3235 => pixel <= "000000";
      when 3236 => pixel <= "000000";
      when 3237 => pixel <= "000000";
      when 3238 => pixel <= "000000";
      when 3239 => pixel <= "000000";
      when 3240 => pixel <= "000000";
      when 3241 => pixel <= "000000";
      when 3242 => pixel <= "000000";
      when 3243 => pixel <= "000000";
      when 3244 => pixel <= "000000";
      when 3245 => pixel <= "000000";
      when 3246 => pixel <= "000000";
      when 3247 => pixel <= "000000";
      when 3248 => pixel <= "000000";
      when 3249 => pixel <= "000000";
      when 3250 => pixel <= "000000";
      when 3251 => pixel <= "000000";
      when 3252 => pixel <= "000000";
      when 3253 => pixel <= "000000";
      when 3254 => pixel <= "000000";
      when 3255 => pixel <= "000000";
      when 3256 => pixel <= "000000";
      when 3257 => pixel <= "000000";
      when 3258 => pixel <= "000000";
      when 3259 => pixel <= "000000";
      when 3260 => pixel <= "000000";
      when 3261 => pixel <= "000000";
      when 3262 => pixel <= "000000";
      when 3263 => pixel <= "000000";
      when 3264 => pixel <= "000000";
      when 3265 => pixel <= "000000";
      when 3266 => pixel <= "000000";
      when 3267 => pixel <= "000000";
      when 3268 => pixel <= "000000";
      when 3269 => pixel <= "000000";
      when 3270 => pixel <= "000000";
      when 3271 => pixel <= "000000";
      when 3272 => pixel <= "000000";
      when 3273 => pixel <= "000000";
      when 3274 => pixel <= "000000";
      when 3275 => pixel <= "000000";
      when 3276 => pixel <= "000000";
      when 3277 => pixel <= "000000";
      when 3278 => pixel <= "000000";
      when 3279 => pixel <= "000000";
      when 3280 => pixel <= "000000";
      when 3281 => pixel <= "000000";
      when 3282 => pixel <= "000000";
      when 3283 => pixel <= "000000";
      when 3284 => pixel <= "000000";
      when 3285 => pixel <= "000000";
      when 3286 => pixel <= "000000";
      when 3287 => pixel <= "000000";
      when 3288 => pixel <= "000000";
      when 3289 => pixel <= "000000";
      when 3290 => pixel <= "000000";
      when 3291 => pixel <= "000000";
      when 3292 => pixel <= "000000";
      when 3293 => pixel <= "000000";
      when 3294 => pixel <= "000000";
      when 3295 => pixel <= "000000";
      when 3296 => pixel <= "000000";
      when 3297 => pixel <= "000000";
      when 3298 => pixel <= "000000";
      when 3299 => pixel <= "000000";
      when 3300 => pixel <= "000000";
      when 3301 => pixel <= "000000";
      when 3302 => pixel <= "000000";
      when 3303 => pixel <= "000000";
      when 3304 => pixel <= "000000";
      when 3305 => pixel <= "000000";
      when 3306 => pixel <= "000000";
      when 3307 => pixel <= "000000";
      when 3308 => pixel <= "000000";
      when 3309 => pixel <= "000000";
      when 3310 => pixel <= "000000";
      when 3311 => pixel <= "000000";
      when 3312 => pixel <= "000000";
      when 3313 => pixel <= "000000";
      when 3314 => pixel <= "000000";
      when 3315 => pixel <= "000000";
      when 3316 => pixel <= "000000";
      when 3317 => pixel <= "000000";
      when 3318 => pixel <= "000000";
      when 3319 => pixel <= "000000";
      when 3320 => pixel <= "000000";
      when 3321 => pixel <= "000000";
      when 3322 => pixel <= "000000";
      when 3323 => pixel <= "000000";
      when 3324 => pixel <= "000000";
      when 3325 => pixel <= "000000";
      when 3326 => pixel <= "000000";
      when 3327 => pixel <= "000000";
      when 3328 => pixel <= "000000";
      when 3329 => pixel <= "000000";
      when 3330 => pixel <= "000000";
      when 3331 => pixel <= "000000";
      when 3332 => pixel <= "000000";
      when 3333 => pixel <= "000000";
      when 3334 => pixel <= "000000";
      when 3335 => pixel <= "000000";
      when 3336 => pixel <= "000000";
      when 3337 => pixel <= "000000";
      when 3338 => pixel <= "000000";
      when 3339 => pixel <= "000000";
      when 3340 => pixel <= "000000";
      when 3341 => pixel <= "000000";
      when 3342 => pixel <= "000000";
      when 3343 => pixel <= "000000";
      when 3344 => pixel <= "000000";
      when 3345 => pixel <= "000000";
      when 3346 => pixel <= "000000";
      when 3347 => pixel <= "000000";
      when 3348 => pixel <= "000000";
      when 3349 => pixel <= "000000";
      when 3350 => pixel <= "000000";
      when 3351 => pixel <= "000000";
      when 3352 => pixel <= "000000";
      when 3353 => pixel <= "000000";
      when 3354 => pixel <= "000000";
      when 3355 => pixel <= "000000";
      when 3356 => pixel <= "000000";
      when 3357 => pixel <= "000000";
      when 3358 => pixel <= "000000";
      when 3359 => pixel <= "000000";
      when 3360 => pixel <= "000000";
      when 3361 => pixel <= "000000";
      when 3362 => pixel <= "000000";
      when 3363 => pixel <= "000000";
      when 3364 => pixel <= "000000";
      when 3365 => pixel <= "000000";
      when 3366 => pixel <= "000000";
      when 3367 => pixel <= "000000";
      when 3368 => pixel <= "000000";
      when 3369 => pixel <= "000000";
      when 3370 => pixel <= "000000";
      when 3371 => pixel <= "000000";
      when 3372 => pixel <= "000000";
      when 3373 => pixel <= "000000";
      when 3374 => pixel <= "000000";
      when 3375 => pixel <= "000000";
      when 3376 => pixel <= "000000";
      when 3377 => pixel <= "000000";
      when 3378 => pixel <= "000000";
      when 3379 => pixel <= "000000";
      when 3380 => pixel <= "000000";
      when 3381 => pixel <= "000000";
      when 3382 => pixel <= "000000";
      when 3383 => pixel <= "000000";
      when 3384 => pixel <= "000000";
      when 3385 => pixel <= "000000";
      when 3386 => pixel <= "000000";
      when 3387 => pixel <= "000000";
      when 3388 => pixel <= "000000";
      when 3389 => pixel <= "000000";
      when 3390 => pixel <= "000000";
      when 3391 => pixel <= "000000";
      when 3392 => pixel <= "000000";
      when 3393 => pixel <= "000000";
      when 3394 => pixel <= "000000";
      when 3395 => pixel <= "000000";
      when 3396 => pixel <= "000000";
      when 3397 => pixel <= "000000";
      when 3398 => pixel <= "000000";
      when 3399 => pixel <= "000000";
      when 3400 => pixel <= "000000";
      when 3401 => pixel <= "000000";
      when 3402 => pixel <= "000000";
      when 3403 => pixel <= "000000";
      when 3404 => pixel <= "000000";
      when 3405 => pixel <= "000000";
      when 3406 => pixel <= "000000";
      when 3407 => pixel <= "000000";
      when 3408 => pixel <= "000000";
      when 3409 => pixel <= "000000";
      when 3410 => pixel <= "000000";
      when 3411 => pixel <= "000000";
      when 3412 => pixel <= "000000";
      when 3413 => pixel <= "000000";
      when 3414 => pixel <= "000000";
      when 3415 => pixel <= "000000";
      when 3416 => pixel <= "000000";
      when 3417 => pixel <= "000000";
      when 3418 => pixel <= "000000";
      when 3419 => pixel <= "000000";
      when 3420 => pixel <= "000000";
      when 3421 => pixel <= "000000";
      when 3422 => pixel <= "000000";
      when 3423 => pixel <= "000000";
      when 3424 => pixel <= "000000";
      when 3425 => pixel <= "000000";
      when 3426 => pixel <= "000000";
      when 3427 => pixel <= "000000";
      when 3428 => pixel <= "000000";
      when 3429 => pixel <= "000000";
      when 3430 => pixel <= "000000";
      when 3431 => pixel <= "000000";
      when 3432 => pixel <= "000000";
      when 3433 => pixel <= "000000";
      when 3434 => pixel <= "000000";
      when 3435 => pixel <= "000000";
      when 3436 => pixel <= "000000";
      when 3437 => pixel <= "000000";
      when 3438 => pixel <= "000000";
      when 3439 => pixel <= "000000";
      when 3440 => pixel <= "000000";
      when 3441 => pixel <= "000000";
      when 3442 => pixel <= "000000";
      when 3443 => pixel <= "000000";
      when 3444 => pixel <= "000000";
      when 3445 => pixel <= "000000";
      when 3446 => pixel <= "000000";
      when 3447 => pixel <= "000000";
      when 3448 => pixel <= "000000";
      when 3449 => pixel <= "000000";
      when 3450 => pixel <= "000000";
      when 3451 => pixel <= "000000";
      when 3452 => pixel <= "000000";
      when 3453 => pixel <= "000000";
      when 3454 => pixel <= "000000";
      when 3455 => pixel <= "000000";
      when 3456 => pixel <= "000000";
      when 3457 => pixel <= "000000";
      when 3458 => pixel <= "000000";
      when 3459 => pixel <= "000000";
      when 3460 => pixel <= "000000";
      when 3461 => pixel <= "000000";
      when 3462 => pixel <= "000000";
      when 3463 => pixel <= "000000";
      when 3464 => pixel <= "000000";
      when 3465 => pixel <= "000000";
      when 3466 => pixel <= "000000";
      when 3467 => pixel <= "000000";
      when 3468 => pixel <= "000000";
      when 3469 => pixel <= "000000";
      when 3470 => pixel <= "000000";
      when 3471 => pixel <= "000000";
      when 3472 => pixel <= "000000";
      when 3473 => pixel <= "000000";
      when 3474 => pixel <= "000000";
      when 3475 => pixel <= "000000";
      when 3476 => pixel <= "000000";
      when 3477 => pixel <= "000000";
      when 3478 => pixel <= "000000";
      when 3479 => pixel <= "000000";
      when 3480 => pixel <= "000000";
      when 3481 => pixel <= "000000";
      when 3482 => pixel <= "000000";
      when 3483 => pixel <= "000000";
      when 3484 => pixel <= "000000";
      when 3485 => pixel <= "000000";
      when 3486 => pixel <= "000000";
      when 3487 => pixel <= "000000";
      when 3488 => pixel <= "000000";
      when 3489 => pixel <= "000000";
      when 3490 => pixel <= "000000";
      when 3491 => pixel <= "000000";
      when 3492 => pixel <= "000000";
      when 3493 => pixel <= "000000";
      when 3494 => pixel <= "000000";
      when 3495 => pixel <= "000000";
      when 3496 => pixel <= "000000";
      when 3497 => pixel <= "000000";
      when 3498 => pixel <= "000000";
      when 3499 => pixel <= "000000";
      when 3500 => pixel <= "000000";
      when 3501 => pixel <= "000000";
      when 3502 => pixel <= "000000";
      when 3503 => pixel <= "000000";
      when 3504 => pixel <= "000000";
      when 3505 => pixel <= "000000";
      when 3506 => pixel <= "000000";
      when 3507 => pixel <= "000000";
      when 3508 => pixel <= "000000";
      when 3509 => pixel <= "000000";
      when 3510 => pixel <= "000000";
      when 3511 => pixel <= "000000";
      when 3512 => pixel <= "000000";
      when 3513 => pixel <= "000000";
      when 3514 => pixel <= "000000";
      when 3515 => pixel <= "000000";
      when 3516 => pixel <= "000000";
      when 3517 => pixel <= "000000";
      when 3518 => pixel <= "000000";
      when 3519 => pixel <= "000000";
      when 3520 => pixel <= "000000";
      when 3521 => pixel <= "000000";
      when 3522 => pixel <= "000000";
      when 3523 => pixel <= "000000";
      when 3524 => pixel <= "000000";
      when 3525 => pixel <= "000000";
      when 3526 => pixel <= "000000";
      when 3527 => pixel <= "000000";
      when 3528 => pixel <= "000000";
      when 3529 => pixel <= "000000";
      when 3530 => pixel <= "000000";
      when 3531 => pixel <= "000000";
      when 3532 => pixel <= "000000";
      when 3533 => pixel <= "000000";
      when 3534 => pixel <= "000000";
      when 3535 => pixel <= "000000";
      when 3536 => pixel <= "000000";
      when 3537 => pixel <= "000000";
      when 3538 => pixel <= "000000";
      when 3539 => pixel <= "000000";
      when 3540 => pixel <= "000000";
      when 3541 => pixel <= "000000";
      when 3542 => pixel <= "000000";
      when 3543 => pixel <= "000000";
      when 3544 => pixel <= "000000";
      when 3545 => pixel <= "000000";
      when 3546 => pixel <= "000000";
      when 3547 => pixel <= "000000";
      when 3548 => pixel <= "000000";
      when 3549 => pixel <= "000000";
      when 3550 => pixel <= "000000";
      when 3551 => pixel <= "000000";
      when 3552 => pixel <= "000000";
      when 3553 => pixel <= "000000";
      when 3554 => pixel <= "000000";
      when 3555 => pixel <= "000000";
      when 3556 => pixel <= "000000";
      when 3557 => pixel <= "000000";
      when 3558 => pixel <= "000000";
      when 3559 => pixel <= "000000";
      when 3560 => pixel <= "000000";
      when 3561 => pixel <= "000000";
      when 3562 => pixel <= "000000";
      when 3563 => pixel <= "000000";
      when 3564 => pixel <= "000000";
      when 3565 => pixel <= "000000";
      when 3566 => pixel <= "000000";
      when 3567 => pixel <= "000000";
      when 3568 => pixel <= "000000";
      when 3569 => pixel <= "000000";
      when 3570 => pixel <= "000000";
      when 3571 => pixel <= "000000";
      when 3572 => pixel <= "000000";
      when 3573 => pixel <= "000000";
      when 3574 => pixel <= "000000";
      when 3575 => pixel <= "000000";
      when 3576 => pixel <= "000000";
      when 3577 => pixel <= "000000";
      when 3578 => pixel <= "000000";
      when 3579 => pixel <= "000000";
      when 3580 => pixel <= "000000";
      when 3581 => pixel <= "000000";
      when 3582 => pixel <= "000000";
      when 3583 => pixel <= "000000";
      when 3584 => pixel <= "000000";
      when 3585 => pixel <= "000000";
      when 3586 => pixel <= "000000";
      when 3587 => pixel <= "000000";
      when 3588 => pixel <= "000000";
      when 3589 => pixel <= "000000";
      when 3590 => pixel <= "000000";
      when 3591 => pixel <= "000000";
      when 3592 => pixel <= "000000";
      when 3593 => pixel <= "000000";
      when 3594 => pixel <= "000000";
      when 3595 => pixel <= "000000";
      when 3596 => pixel <= "000000";
      when 3597 => pixel <= "000000";
      when 3598 => pixel <= "000000";
      when 3599 => pixel <= "000000";
      when 3600 => pixel <= "000000";
      when 3601 => pixel <= "000000";
      when 3602 => pixel <= "000000";
      when 3603 => pixel <= "000000";
      when 3604 => pixel <= "000000";
      when 3605 => pixel <= "000000";
      when 3606 => pixel <= "000000";
      when 3607 => pixel <= "000000";
      when 3608 => pixel <= "000000";
      when 3609 => pixel <= "000000";
      when 3610 => pixel <= "000000";
      when 3611 => pixel <= "000000";
      when 3612 => pixel <= "000000";
      when 3613 => pixel <= "000000";
      when 3614 => pixel <= "000000";
      when 3615 => pixel <= "000000";
      when 3616 => pixel <= "000000";
      when 3617 => pixel <= "000000";
      when 3618 => pixel <= "000000";
      when 3619 => pixel <= "000000";
      when 3620 => pixel <= "000000";
      when 3621 => pixel <= "000000";
      when 3622 => pixel <= "000000";
      when 3623 => pixel <= "000000";
      when 3624 => pixel <= "000000";
      when 3625 => pixel <= "000000";
      when 3626 => pixel <= "000000";
      when 3627 => pixel <= "000000";
      when 3628 => pixel <= "000000";
      when 3629 => pixel <= "000000";
      when 3630 => pixel <= "000000";
      when 3631 => pixel <= "000000";
      when 3632 => pixel <= "000000";
      when 3633 => pixel <= "000000";
      when 3634 => pixel <= "000000";
      when 3635 => pixel <= "000000";
      when 3636 => pixel <= "000000";
      when 3637 => pixel <= "000000";
      when 3638 => pixel <= "000000";
      when 3639 => pixel <= "000000";
      when 3640 => pixel <= "000000";
      when 3641 => pixel <= "000000";
      when 3642 => pixel <= "000000";
      when 3643 => pixel <= "000000";
      when 3644 => pixel <= "000000";
      when 3645 => pixel <= "000000";
      when 3646 => pixel <= "000000";
      when 3647 => pixel <= "000000";
      when 3648 => pixel <= "000000";
      when 3649 => pixel <= "000000";
      when 3650 => pixel <= "000000";
      when 3651 => pixel <= "000000";
      when 3652 => pixel <= "000000";
      when 3653 => pixel <= "000000";
      when 3654 => pixel <= "000000";
      when 3655 => pixel <= "000000";
      when 3656 => pixel <= "000000";
      when 3657 => pixel <= "000000";
      when 3658 => pixel <= "000000";
      when 3659 => pixel <= "000000";
      when 3660 => pixel <= "000000";
      when 3661 => pixel <= "000000";
      when 3662 => pixel <= "000000";
      when 3663 => pixel <= "000000";
      when 3664 => pixel <= "000000";
      when 3665 => pixel <= "000000";
      when 3666 => pixel <= "000000";
      when 3667 => pixel <= "000000";
      when 3668 => pixel <= "000000";
      when 3669 => pixel <= "000000";
      when 3670 => pixel <= "000000";
      when 3671 => pixel <= "000000";
      when 3672 => pixel <= "000000";
      when 3673 => pixel <= "000000";
      when 3674 => pixel <= "000000";
      when 3675 => pixel <= "000000";
      when 3676 => pixel <= "000000";
      when 3677 => pixel <= "000000";
      when 3678 => pixel <= "000000";
      when 3679 => pixel <= "000000";
      when 3680 => pixel <= "000000";
      when 3681 => pixel <= "000000";
      when 3682 => pixel <= "000000";
      when 3683 => pixel <= "000000";
      when 3684 => pixel <= "000000";
      when 3685 => pixel <= "000000";
      when 3686 => pixel <= "000000";
      when 3687 => pixel <= "000000";
      when 3688 => pixel <= "000000";
      when 3689 => pixel <= "000000";
      when 3690 => pixel <= "000000";
      when 3691 => pixel <= "000000";
      when 3692 => pixel <= "000000";
      when 3693 => pixel <= "000000";
      when 3694 => pixel <= "000000";
      when 3695 => pixel <= "000000";
      when 3696 => pixel <= "000000";
      when 3697 => pixel <= "000000";
      when 3698 => pixel <= "000000";
      when 3699 => pixel <= "000000";
      when 3700 => pixel <= "000000";
      when 3701 => pixel <= "000000";
      when 3702 => pixel <= "000000";
      when 3703 => pixel <= "000000";
      when 3704 => pixel <= "000000";
      when 3705 => pixel <= "000000";
      when 3706 => pixel <= "000000";
      when 3707 => pixel <= "000000";
      when 3708 => pixel <= "000000";
      when 3709 => pixel <= "000000";
      when 3710 => pixel <= "000000";
      when 3711 => pixel <= "000000";
      when 3712 => pixel <= "000000";
      when 3713 => pixel <= "000000";
      when 3714 => pixel <= "000000";
      when 3715 => pixel <= "000000";
      when 3716 => pixel <= "000000";
      when 3717 => pixel <= "000000";
      when 3718 => pixel <= "000000";
      when 3719 => pixel <= "000000";
      when 3720 => pixel <= "000000";
      when 3721 => pixel <= "000000";
      when 3722 => pixel <= "000000";
      when 3723 => pixel <= "000000";
      when 3724 => pixel <= "000000";
      when 3725 => pixel <= "000000";
      when 3726 => pixel <= "000000";
      when 3727 => pixel <= "000000";
      when 3728 => pixel <= "000000";
      when 3729 => pixel <= "000000";
      when 3730 => pixel <= "000000";
      when 3731 => pixel <= "000000";
      when 3732 => pixel <= "000000";
      when 3733 => pixel <= "000000";
      when 3734 => pixel <= "000000";
      when 3735 => pixel <= "000000";
      when 3736 => pixel <= "000000";
      when 3737 => pixel <= "000000";
      when 3738 => pixel <= "000000";
      when 3739 => pixel <= "000000";
      when 3740 => pixel <= "000000";
      when 3741 => pixel <= "000000";
      when 3742 => pixel <= "000000";
      when 3743 => pixel <= "000000";
      when 3744 => pixel <= "000000";
      when 3745 => pixel <= "000000";
      when 3746 => pixel <= "000000";
      when 3747 => pixel <= "000000";
      when 3748 => pixel <= "000000";
      when 3749 => pixel <= "000000";
      when 3750 => pixel <= "000000";
      when 3751 => pixel <= "000000";
      when 3752 => pixel <= "000000";
      when 3753 => pixel <= "000000";
      when 3754 => pixel <= "000000";
      when 3755 => pixel <= "000000";
      when 3756 => pixel <= "000000";
      when 3757 => pixel <= "000000";
      when 3758 => pixel <= "000000";
      when 3759 => pixel <= "000000";
      when 3760 => pixel <= "000000";
      when 3761 => pixel <= "000000";
      when 3762 => pixel <= "000000";
      when 3763 => pixel <= "000000";
      when 3764 => pixel <= "000000";
      when 3765 => pixel <= "000000";
      when 3766 => pixel <= "000000";
      when 3767 => pixel <= "000000";
      when 3768 => pixel <= "000000";
      when 3769 => pixel <= "000000";
      when 3770 => pixel <= "000000";
      when 3771 => pixel <= "000000";
      when 3772 => pixel <= "000000";
      when 3773 => pixel <= "000000";
      when 3774 => pixel <= "000000";
      when 3775 => pixel <= "000000";
      when 3776 => pixel <= "000000";
      when 3777 => pixel <= "000000";
      when 3778 => pixel <= "000000";
      when 3779 => pixel <= "000000";
      when 3780 => pixel <= "000000";
      when 3781 => pixel <= "000000";
      when 3782 => pixel <= "000000";
      when 3783 => pixel <= "000000";
      when 3784 => pixel <= "000000";
      when 3785 => pixel <= "000000";
      when 3786 => pixel <= "000000";
      when 3787 => pixel <= "000000";
      when 3788 => pixel <= "000000";
      when 3789 => pixel <= "000000";
      when 3790 => pixel <= "000000";
      when 3791 => pixel <= "000000";
      when 3792 => pixel <= "000000";
      when 3793 => pixel <= "000000";
      when 3794 => pixel <= "000000";
      when 3795 => pixel <= "000000";
      when 3796 => pixel <= "000000";
      when 3797 => pixel <= "000000";
      when 3798 => pixel <= "000000";
      when 3799 => pixel <= "000000";
      when 3800 => pixel <= "000000";
      when 3801 => pixel <= "000000";
      when 3802 => pixel <= "000000";
      when 3803 => pixel <= "000000";
      when 3804 => pixel <= "000000";
      when 3805 => pixel <= "000000";
      when 3806 => pixel <= "000000";
      when 3807 => pixel <= "000000";
      when 3808 => pixel <= "000000";
      when 3809 => pixel <= "000000";
      when 3810 => pixel <= "000000";
      when 3811 => pixel <= "000000";
      when 3812 => pixel <= "000000";
      when 3813 => pixel <= "000000";
      when 3814 => pixel <= "000000";
      when 3815 => pixel <= "000000";
      when 3816 => pixel <= "000000";
      when 3817 => pixel <= "000000";
      when 3818 => pixel <= "000000";
      when 3819 => pixel <= "000000";
      when 3820 => pixel <= "000000";
      when 3821 => pixel <= "000000";
      when 3822 => pixel <= "000000";
      when 3823 => pixel <= "000000";
      when 3824 => pixel <= "000000";
      when 3825 => pixel <= "000000";
      when 3826 => pixel <= "000000";
      when 3827 => pixel <= "000000";
      when 3828 => pixel <= "000000";
      when 3829 => pixel <= "000000";
      when 3830 => pixel <= "000000";
      when 3831 => pixel <= "000000";
      when 3832 => pixel <= "000000";
      when 3833 => pixel <= "000000";
      when 3834 => pixel <= "000000";
      when 3835 => pixel <= "000000";
      when 3836 => pixel <= "000000";
      when 3837 => pixel <= "000000";
      when 3838 => pixel <= "000000";
      when 3839 => pixel <= "000000";
      when 3840 => pixel <= "000000";
      when 3841 => pixel <= "000000";
      when 3842 => pixel <= "000000";
      when 3843 => pixel <= "000000";
      when 3844 => pixel <= "000000";
      when 3845 => pixel <= "000000";
      when 3846 => pixel <= "000000";
      when 3847 => pixel <= "000000";
      when 3848 => pixel <= "000000";
      when 3849 => pixel <= "000000";
      when 3850 => pixel <= "000000";
      when 3851 => pixel <= "000000";
      when 3852 => pixel <= "000000";
      when 3853 => pixel <= "000000";
      when 3854 => pixel <= "000000";
      when 3855 => pixel <= "000000";
      when 3856 => pixel <= "000000";
      when 3857 => pixel <= "000000";
      when 3858 => pixel <= "000000";
      when 3859 => pixel <= "000000";
      when 3860 => pixel <= "000000";
      when 3861 => pixel <= "000000";
      when 3862 => pixel <= "000000";
      when 3863 => pixel <= "000000";
      when 3864 => pixel <= "000000";
      when 3865 => pixel <= "000000";
      when 3866 => pixel <= "000000";
      when 3867 => pixel <= "000000";
      when 3868 => pixel <= "000000";
      when 3869 => pixel <= "000000";
      when 3870 => pixel <= "000000";
      when 3871 => pixel <= "000000";
      when 3872 => pixel <= "000000";
      when 3873 => pixel <= "000000";
      when 3874 => pixel <= "000000";
      when 3875 => pixel <= "000000";
      when 3876 => pixel <= "000000";
      when 3877 => pixel <= "000000";
      when 3878 => pixel <= "000000";
      when 3879 => pixel <= "000000";
      when 3880 => pixel <= "000000";
      when 3881 => pixel <= "000000";
      when 3882 => pixel <= "000000";
      when 3883 => pixel <= "000000";
      when 3884 => pixel <= "000000";
      when 3885 => pixel <= "000000";
      when 3886 => pixel <= "000000";
      when 3887 => pixel <= "000000";
      when 3888 => pixel <= "000000";
      when 3889 => pixel <= "000000";
      when 3890 => pixel <= "000000";
      when 3891 => pixel <= "000000";
      when 3892 => pixel <= "000000";
      when 3893 => pixel <= "000000";
      when 3894 => pixel <= "000000";
      when 3895 => pixel <= "000000";
      when 3896 => pixel <= "000000";
      when 3897 => pixel <= "000000";
      when 3898 => pixel <= "000000";
      when 3899 => pixel <= "000000";
      when 3900 => pixel <= "000000";
      when 3901 => pixel <= "000000";
      when 3902 => pixel <= "000000";
      when 3903 => pixel <= "000000";
      when 3904 => pixel <= "000000";
      when 3905 => pixel <= "000000";
      when 3906 => pixel <= "000000";
      when 3907 => pixel <= "000000";
      when 3908 => pixel <= "000000";
      when 3909 => pixel <= "000000";
      when 3910 => pixel <= "000000";
      when 3911 => pixel <= "000000";
      when 3912 => pixel <= "000000";
      when 3913 => pixel <= "000000";
      when 3914 => pixel <= "000000";
      when 3915 => pixel <= "000000";
      when 3916 => pixel <= "000000";
      when 3917 => pixel <= "000000";
      when 3918 => pixel <= "000000";
      when 3919 => pixel <= "000000";
      when 3920 => pixel <= "000000";
      when 3921 => pixel <= "000000";
      when 3922 => pixel <= "000000";
      when 3923 => pixel <= "000000";
      when 3924 => pixel <= "000000";
      when 3925 => pixel <= "000000";
      when 3926 => pixel <= "000000";
      when 3927 => pixel <= "000000";
      when 3928 => pixel <= "000000";
      when 3929 => pixel <= "000000";
      when 3930 => pixel <= "000000";
      when 3931 => pixel <= "000000";
      when 3932 => pixel <= "000000";
      when 3933 => pixel <= "000000";
      when 3934 => pixel <= "000000";
      when 3935 => pixel <= "000000";
      when 3936 => pixel <= "000000";
      when 3937 => pixel <= "000000";
      when 3938 => pixel <= "000000";
      when 3939 => pixel <= "000000";
      when 3940 => pixel <= "000000";
      when 3941 => pixel <= "000000";
      when 3942 => pixel <= "000000";
      when 3943 => pixel <= "000000";
      when 3944 => pixel <= "000000";
      when 3945 => pixel <= "000000";
      when 3946 => pixel <= "000000";
      when 3947 => pixel <= "000000";
      when 3948 => pixel <= "000000";
      when 3949 => pixel <= "000000";
      when 3950 => pixel <= "000000";
      when 3951 => pixel <= "000000";
      when 3952 => pixel <= "000000";
      when 3953 => pixel <= "000000";
      when 3954 => pixel <= "000000";
      when 3955 => pixel <= "000000";
      when 3956 => pixel <= "000000";
      when 3957 => pixel <= "000000";
      when 3958 => pixel <= "000000";
      when 3959 => pixel <= "000000";
      when 3960 => pixel <= "000000";
      when 3961 => pixel <= "000000";
      when 3962 => pixel <= "000000";
      when 3963 => pixel <= "000000";
      when 3964 => pixel <= "000000";
      when 3965 => pixel <= "000000";
      when 3966 => pixel <= "000000";
      when 3967 => pixel <= "000000";
      when 3968 => pixel <= "000000";
      when 3969 => pixel <= "000000";
      when 3970 => pixel <= "000000";
      when 3971 => pixel <= "000000";
      when 3972 => pixel <= "000000";
      when 3973 => pixel <= "000000";
      when 3974 => pixel <= "000000";
      when 3975 => pixel <= "000000";
      when 3976 => pixel <= "000000";
      when 3977 => pixel <= "000000";
      when 3978 => pixel <= "000000";
      when 3979 => pixel <= "000000";
      when 3980 => pixel <= "000000";
      when 3981 => pixel <= "000000";
      when 3982 => pixel <= "000000";
      when 3983 => pixel <= "000000";
      when 3984 => pixel <= "000000";
      when 3985 => pixel <= "000000";
      when 3986 => pixel <= "000000";
      when 3987 => pixel <= "000000";
      when 3988 => pixel <= "000000";
      when 3989 => pixel <= "000000";
      when 3990 => pixel <= "000000";
      when 3991 => pixel <= "000000";
      when 3992 => pixel <= "000000";
      when 3993 => pixel <= "000000";
      when 3994 => pixel <= "000000";
      when 3995 => pixel <= "000000";
      when 3996 => pixel <= "000000";
      when 3997 => pixel <= "000000";
      when 3998 => pixel <= "000000";
      when 3999 => pixel <= "000000";
      when 4000 => pixel <= "000000";
      when 4001 => pixel <= "000000";
      when 4002 => pixel <= "000000";
      when 4003 => pixel <= "000000";
      when 4004 => pixel <= "000000";
      when 4005 => pixel <= "000000";
      when 4006 => pixel <= "000000";
      when 4007 => pixel <= "000000";
      when 4008 => pixel <= "000000";
      when 4009 => pixel <= "000000";
      when 4010 => pixel <= "000000";
      when 4011 => pixel <= "000000";
      when 4012 => pixel <= "000000";
      when 4013 => pixel <= "000000";
      when 4014 => pixel <= "000000";
      when 4015 => pixel <= "000000";
      when 4016 => pixel <= "000000";
      when 4017 => pixel <= "000000";
      when 4018 => pixel <= "000000";
      when 4019 => pixel <= "000000";
      when 4020 => pixel <= "000000";
      when 4021 => pixel <= "000000";
      when 4022 => pixel <= "000000";
      when 4023 => pixel <= "000000";
      when 4024 => pixel <= "000000";
      when 4025 => pixel <= "000000";
      when 4026 => pixel <= "000000";
      when 4027 => pixel <= "000000";
      when 4028 => pixel <= "000000";
      when 4029 => pixel <= "000000";
      when 4030 => pixel <= "000000";
      when 4031 => pixel <= "000000";
      when 4032 => pixel <= "000000";
      when 4033 => pixel <= "000000";
      when 4034 => pixel <= "000000";
      when 4035 => pixel <= "000000";
      when 4036 => pixel <= "000000";
      when 4037 => pixel <= "000000";
      when 4038 => pixel <= "000000";
      when 4039 => pixel <= "000000";
      when 4040 => pixel <= "000000";
      when 4041 => pixel <= "000000";
      when 4042 => pixel <= "000000";
      when 4043 => pixel <= "000000";
      when 4044 => pixel <= "000000";
      when 4045 => pixel <= "000000";
      when 4046 => pixel <= "000000";
      when 4047 => pixel <= "000000";
      when 4048 => pixel <= "000000";
      when 4049 => pixel <= "000000";
      when 4050 => pixel <= "000000";
      when 4051 => pixel <= "000000";
      when 4052 => pixel <= "000000";
      when 4053 => pixel <= "000000";
      when 4054 => pixel <= "000000";
      when 4055 => pixel <= "000000";
      when 4056 => pixel <= "000000";
      when 4057 => pixel <= "000000";
      when 4058 => pixel <= "000000";
      when 4059 => pixel <= "000000";
      when 4060 => pixel <= "000000";
      when 4061 => pixel <= "000000";
      when 4062 => pixel <= "000000";
      when 4063 => pixel <= "000000";
      when 4064 => pixel <= "000000";
      when 4065 => pixel <= "000000";
      when 4066 => pixel <= "000000";
      when 4067 => pixel <= "000000";
      when 4068 => pixel <= "000000";
      when 4069 => pixel <= "000000";
      when 4070 => pixel <= "000000";
      when 4071 => pixel <= "000000";
      when 4072 => pixel <= "000000";
      when 4073 => pixel <= "000000";
      when 4074 => pixel <= "000000";
      when 4075 => pixel <= "000000";
      when 4076 => pixel <= "000000";
      when 4077 => pixel <= "000000";
      when 4078 => pixel <= "000000";
      when 4079 => pixel <= "000000";
      when 4080 => pixel <= "000000";
      when 4081 => pixel <= "000000";
      when 4082 => pixel <= "000000";
      when 4083 => pixel <= "000000";
      when 4084 => pixel <= "000000";
      when 4085 => pixel <= "000000";
      when 4086 => pixel <= "000000";
      when 4087 => pixel <= "000000";
      when 4088 => pixel <= "000000";
      when 4089 => pixel <= "000000";
      when 4090 => pixel <= "000000";
      when 4091 => pixel <= "000000";
      when 4092 => pixel <= "000000";
      when 4093 => pixel <= "000000";
      when 4094 => pixel <= "000000";
      when 4095 => pixel <= "000000";
      when 4096 => pixel <= "000000";
      when 4097 => pixel <= "000000";
      when 4098 => pixel <= "000000";
      when 4099 => pixel <= "000000";
      when 4100 => pixel <= "000000";
      when 4101 => pixel <= "000000";
      when 4102 => pixel <= "000000";
      when 4103 => pixel <= "000000";
      when 4104 => pixel <= "000000";
      when 4105 => pixel <= "000000";
      when 4106 => pixel <= "000000";
      when 4107 => pixel <= "000000";
      when 4108 => pixel <= "000000";
      when 4109 => pixel <= "000000";
      when 4110 => pixel <= "000000";
      when 4111 => pixel <= "000000";
      when 4112 => pixel <= "000000";
      when 4113 => pixel <= "000000";
      when 4114 => pixel <= "000000";
      when 4115 => pixel <= "000000";
      when 4116 => pixel <= "000000";
      when 4117 => pixel <= "000000";
      when 4118 => pixel <= "000000";
      when 4119 => pixel <= "000000";
      when 4120 => pixel <= "000000";
      when 4121 => pixel <= "000000";
      when 4122 => pixel <= "000000";
      when 4123 => pixel <= "000000";
      when 4124 => pixel <= "000000";
      when 4125 => pixel <= "000000";
      when 4126 => pixel <= "000000";
      when 4127 => pixel <= "000000";
      when 4128 => pixel <= "000000";
      when 4129 => pixel <= "000000";
      when 4130 => pixel <= "000000";
      when 4131 => pixel <= "000000";
      when 4132 => pixel <= "000000";
      when 4133 => pixel <= "000000";
      when 4134 => pixel <= "000000";
      when 4135 => pixel <= "000000";
      when 4136 => pixel <= "000000";
      when 4137 => pixel <= "000000";
      when 4138 => pixel <= "000000";
      when 4139 => pixel <= "000000";
      when 4140 => pixel <= "000000";
      when 4141 => pixel <= "000000";
      when 4142 => pixel <= "000000";
      when 4143 => pixel <= "000000";
      when 4144 => pixel <= "000000";
      when 4145 => pixel <= "000000";
      when 4146 => pixel <= "000000";
      when 4147 => pixel <= "000000";
      when 4148 => pixel <= "000000";
      when 4149 => pixel <= "000000";
      when 4150 => pixel <= "000000";
      when 4151 => pixel <= "000000";
      when 4152 => pixel <= "000000";
      when 4153 => pixel <= "000000";
      when 4154 => pixel <= "000000";
      when 4155 => pixel <= "000000";
      when 4156 => pixel <= "000000";
      when 4157 => pixel <= "000000";
      when 4158 => pixel <= "000000";
      when 4159 => pixel <= "000000";
      when 4160 => pixel <= "000000";
      when 4161 => pixel <= "000000";
      when 4162 => pixel <= "000000";
      when 4163 => pixel <= "000000";
      when 4164 => pixel <= "000000";
      when 4165 => pixel <= "000000";
      when 4166 => pixel <= "000000";
      when 4167 => pixel <= "000000";
      when 4168 => pixel <= "000000";
      when 4169 => pixel <= "000000";
      when 4170 => pixel <= "000000";
      when 4171 => pixel <= "000000";
      when 4172 => pixel <= "000000";
      when 4173 => pixel <= "000000";
      when 4174 => pixel <= "000000";
      when 4175 => pixel <= "000000";
      when 4176 => pixel <= "000000";
      when 4177 => pixel <= "000000";
      when 4178 => pixel <= "000000";
      when 4179 => pixel <= "000000";
      when 4180 => pixel <= "000000";
      when 4181 => pixel <= "000000";
      when 4182 => pixel <= "000000";
      when 4183 => pixel <= "000000";
      when 4184 => pixel <= "000000";
      when 4185 => pixel <= "000000";
      when 4186 => pixel <= "000000";
      when 4187 => pixel <= "000000";
      when 4188 => pixel <= "000000";
      when 4189 => pixel <= "000000";
      when 4190 => pixel <= "000000";
      when 4191 => pixel <= "000000";
      when 4192 => pixel <= "000000";
      when 4193 => pixel <= "000000";
      when 4194 => pixel <= "000000";
      when 4195 => pixel <= "000000";
      when 4196 => pixel <= "000000";
      when 4197 => pixel <= "000000";
      when 4198 => pixel <= "000000";
      when 4199 => pixel <= "000000";
      when 4200 => pixel <= "000000";
      when 4201 => pixel <= "000000";
      when 4202 => pixel <= "000000";
      when 4203 => pixel <= "000000";
      when 4204 => pixel <= "000000";
      when 4205 => pixel <= "000000";
      when 4206 => pixel <= "000000";
      when 4207 => pixel <= "000000";
      when 4208 => pixel <= "000000";
      when 4209 => pixel <= "000000";
      when 4210 => pixel <= "000000";
      when 4211 => pixel <= "000000";
      when 4212 => pixel <= "000000";
      when 4213 => pixel <= "000000";
      when 4214 => pixel <= "000000";
      when 4215 => pixel <= "000000";
      when 4216 => pixel <= "000000";
      when 4217 => pixel <= "000000";
      when 4218 => pixel <= "000000";
      when 4219 => pixel <= "000000";
      when 4220 => pixel <= "000000";
      when 4221 => pixel <= "000000";
      when 4222 => pixel <= "000000";
      when 4223 => pixel <= "000000";
      when 4224 => pixel <= "000000";
      when 4225 => pixel <= "000000";
      when 4226 => pixel <= "000000";
      when 4227 => pixel <= "000000";
      when 4228 => pixel <= "000000";
      when 4229 => pixel <= "000000";
      when 4230 => pixel <= "000000";
      when 4231 => pixel <= "000000";
      when 4232 => pixel <= "000000";
      when 4233 => pixel <= "000000";
      when 4234 => pixel <= "000000";
      when 4235 => pixel <= "000000";
      when 4236 => pixel <= "000000";
      when 4237 => pixel <= "000000";
      when 4238 => pixel <= "000000";
      when 4239 => pixel <= "000000";
      when 4240 => pixel <= "000000";
      when 4241 => pixel <= "000000";
      when 4242 => pixel <= "000000";
      when 4243 => pixel <= "000000";
      when 4244 => pixel <= "000000";
      when 4245 => pixel <= "000000";
      when 4246 => pixel <= "000000";
      when 4247 => pixel <= "000000";
      when 4248 => pixel <= "000000";
      when 4249 => pixel <= "000000";
      when 4250 => pixel <= "000000";
      when 4251 => pixel <= "000000";
      when 4252 => pixel <= "000000";
      when 4253 => pixel <= "000000";
      when 4254 => pixel <= "000000";
      when 4255 => pixel <= "000000";
      when 4256 => pixel <= "000000";
      when 4257 => pixel <= "000000";
      when 4258 => pixel <= "000000";
      when 4259 => pixel <= "000000";
      when 4260 => pixel <= "000000";
      when 4261 => pixel <= "000000";
      when 4262 => pixel <= "000000";
      when 4263 => pixel <= "000000";
      when 4264 => pixel <= "000000";
      when 4265 => pixel <= "000000";
      when 4266 => pixel <= "000000";
      when 4267 => pixel <= "000000";
      when 4268 => pixel <= "000000";
      when 4269 => pixel <= "000000";
      when 4270 => pixel <= "000000";
      when 4271 => pixel <= "000000";
      when 4272 => pixel <= "000000";
      when 4273 => pixel <= "000000";
      when 4274 => pixel <= "000000";
      when 4275 => pixel <= "000000";
      when 4276 => pixel <= "000000";
      when 4277 => pixel <= "000000";
      when 4278 => pixel <= "000000";
      when 4279 => pixel <= "000000";
      when 4280 => pixel <= "000000";
      when 4281 => pixel <= "000000";
      when 4282 => pixel <= "000000";
      when 4283 => pixel <= "000000";
      when 4284 => pixel <= "000000";
      when 4285 => pixel <= "000000";
      when 4286 => pixel <= "000000";
      when 4287 => pixel <= "000000";
      when 4288 => pixel <= "000000";
      when 4289 => pixel <= "000000";
      when 4290 => pixel <= "000000";
      when 4291 => pixel <= "000000";
      when 4292 => pixel <= "000000";
      when 4293 => pixel <= "000000";
      when 4294 => pixel <= "000000";
      when 4295 => pixel <= "000000";
      when 4296 => pixel <= "000000";
      when 4297 => pixel <= "000000";
      when 4298 => pixel <= "000000";
      when 4299 => pixel <= "000000";
      when 4300 => pixel <= "000000";
      when 4301 => pixel <= "000000";
      when 4302 => pixel <= "000000";
      when 4303 => pixel <= "000000";
      when 4304 => pixel <= "000000";
      when 4305 => pixel <= "000000";
      when 4306 => pixel <= "000000";
      when 4307 => pixel <= "000000";
      when 4308 => pixel <= "000000";
      when 4309 => pixel <= "000000";
      when 4310 => pixel <= "000000";
      when 4311 => pixel <= "000000";
      when 4312 => pixel <= "000000";
      when 4313 => pixel <= "000000";
      when 4314 => pixel <= "000000";
      when 4315 => pixel <= "000000";
      when 4316 => pixel <= "000000";
      when 4317 => pixel <= "000000";
      when 4318 => pixel <= "000000";
      when 4319 => pixel <= "000000";
      when 4320 => pixel <= "000000";
      when 4321 => pixel <= "000000";
      when 4322 => pixel <= "000000";
      when 4323 => pixel <= "000000";
      when 4324 => pixel <= "000000";
      when 4325 => pixel <= "000000";
      when 4326 => pixel <= "000000";
      when 4327 => pixel <= "000000";
      when 4328 => pixel <= "000000";
      when 4329 => pixel <= "000000";
      when 4330 => pixel <= "000000";
      when 4331 => pixel <= "000000";
      when 4332 => pixel <= "000000";
      when 4333 => pixel <= "000000";
      when 4334 => pixel <= "000000";
      when 4335 => pixel <= "000000";
      when 4336 => pixel <= "000000";
      when 4337 => pixel <= "000000";
      when 4338 => pixel <= "000000";
      when 4339 => pixel <= "000000";
      when 4340 => pixel <= "000000";
      when 4341 => pixel <= "000000";
      when 4342 => pixel <= "000000";
      when 4343 => pixel <= "000000";
      when 4344 => pixel <= "000000";
      when 4345 => pixel <= "000000";
      when 4346 => pixel <= "000000";
      when 4347 => pixel <= "000000";
      when 4348 => pixel <= "000000";
      when 4349 => pixel <= "000000";
      when 4350 => pixel <= "000000";
      when 4351 => pixel <= "000000";
      when 4352 => pixel <= "000000";
      when 4353 => pixel <= "000000";
      when 4354 => pixel <= "000000";
      when 4355 => pixel <= "000000";
      when 4356 => pixel <= "000000";
      when 4357 => pixel <= "000000";
      when 4358 => pixel <= "000000";
      when 4359 => pixel <= "000000";
      when 4360 => pixel <= "000000";
      when 4361 => pixel <= "000000";
      when 4362 => pixel <= "000000";
      when 4363 => pixel <= "000000";
      when 4364 => pixel <= "000000";
      when 4365 => pixel <= "000000";
      when 4366 => pixel <= "000000";
      when 4367 => pixel <= "000000";
      when 4368 => pixel <= "000000";
      when 4369 => pixel <= "000000";
      when 4370 => pixel <= "000000";
      when 4371 => pixel <= "000000";
      when 4372 => pixel <= "000000";
      when 4373 => pixel <= "000000";
      when 4374 => pixel <= "000000";
      when 4375 => pixel <= "000000";
      when 4376 => pixel <= "000000";
      when 4377 => pixel <= "000000";
      when 4378 => pixel <= "000000";
      when 4379 => pixel <= "000000";
      when 4380 => pixel <= "000000";
      when 4381 => pixel <= "000000";
      when 4382 => pixel <= "000000";
      when 4383 => pixel <= "000000";
      when 4384 => pixel <= "000000";
      when 4385 => pixel <= "000000";
      when 4386 => pixel <= "000000";
      when 4387 => pixel <= "000000";
      when 4388 => pixel <= "000000";
      when 4389 => pixel <= "000000";
      when 4390 => pixel <= "000000";
      when 4391 => pixel <= "000000";
      when 4392 => pixel <= "000000";
      when 4393 => pixel <= "000000";
      when 4394 => pixel <= "000000";
      when 4395 => pixel <= "000000";
      when 4396 => pixel <= "000000";
      when 4397 => pixel <= "000000";
      when 4398 => pixel <= "000000";
      when 4399 => pixel <= "000000";
      when 4400 => pixel <= "000000";
      when 4401 => pixel <= "000000";
      when 4402 => pixel <= "000000";
      when 4403 => pixel <= "000000";
      when 4404 => pixel <= "000000";
      when 4405 => pixel <= "000000";
      when 4406 => pixel <= "000000";
      when 4407 => pixel <= "000000";
      when 4408 => pixel <= "000000";
      when 4409 => pixel <= "000000";
      when 4410 => pixel <= "000000";
      when 4411 => pixel <= "000000";
      when 4412 => pixel <= "000000";
      when 4413 => pixel <= "000000";
      when 4414 => pixel <= "000000";
      when 4415 => pixel <= "000000";
      when 4416 => pixel <= "000000";
      when 4417 => pixel <= "000000";
      when 4418 => pixel <= "000000";
      when 4419 => pixel <= "000000";
      when 4420 => pixel <= "000000";
      when 4421 => pixel <= "000000";
      when 4422 => pixel <= "000000";
      when 4423 => pixel <= "000000";
      when 4424 => pixel <= "000000";
      when 4425 => pixel <= "000000";
      when 4426 => pixel <= "000000";
      when 4427 => pixel <= "000000";
      when 4428 => pixel <= "000000";
      when 4429 => pixel <= "000000";
      when 4430 => pixel <= "000000";
      when 4431 => pixel <= "000000";
      when 4432 => pixel <= "000000";
      when 4433 => pixel <= "000000";
      when 4434 => pixel <= "000000";
      when 4435 => pixel <= "000000";
      when 4436 => pixel <= "000000";
      when 4437 => pixel <= "000000";
      when 4438 => pixel <= "000000";
      when 4439 => pixel <= "000000";
      when 4440 => pixel <= "000000";
      when 4441 => pixel <= "000000";
      when 4442 => pixel <= "000000";
      when 4443 => pixel <= "000000";
      when 4444 => pixel <= "000000";
      when 4445 => pixel <= "000000";
      when 4446 => pixel <= "000000";
      when 4447 => pixel <= "000000";
      when 4448 => pixel <= "000000";
      when 4449 => pixel <= "000000";
      when 4450 => pixel <= "000000";
      when 4451 => pixel <= "000000";
      when 4452 => pixel <= "000000";
      when 4453 => pixel <= "000000";
      when 4454 => pixel <= "000000";
      when 4455 => pixel <= "000000";
      when 4456 => pixel <= "000000";
      when 4457 => pixel <= "000000";
      when 4458 => pixel <= "000000";
      when 4459 => pixel <= "000000";
      when 4460 => pixel <= "000000";
      when 4461 => pixel <= "000000";
      when 4462 => pixel <= "000000";
      when 4463 => pixel <= "000000";
      when 4464 => pixel <= "000000";
      when 4465 => pixel <= "000000";
      when 4466 => pixel <= "000000";
      when 4467 => pixel <= "000000";
      when 4468 => pixel <= "000000";
      when 4469 => pixel <= "000000";
      when 4470 => pixel <= "000000";
      when 4471 => pixel <= "000000";
      when 4472 => pixel <= "000000";
      when 4473 => pixel <= "000000";
      when 4474 => pixel <= "000000";
      when 4475 => pixel <= "000000";
      when 4476 => pixel <= "000000";
      when 4477 => pixel <= "000000";
      when 4478 => pixel <= "000000";
      when 4479 => pixel <= "000000";
      when 4480 => pixel <= "000000";
      when 4481 => pixel <= "000000";
      when 4482 => pixel <= "000000";
      when 4483 => pixel <= "000000";
      when 4484 => pixel <= "000000";
      when 4485 => pixel <= "000000";
      when 4486 => pixel <= "000000";
      when 4487 => pixel <= "000000";
      when 4488 => pixel <= "000000";
      when 4489 => pixel <= "000000";
      when 4490 => pixel <= "000000";
      when 4491 => pixel <= "000000";
      when 4492 => pixel <= "000000";
      when 4493 => pixel <= "000000";
      when 4494 => pixel <= "000000";
      when 4495 => pixel <= "000000";
      when 4496 => pixel <= "000000";
      when 4497 => pixel <= "000000";
      when 4498 => pixel <= "000000";
      when 4499 => pixel <= "000000";
      when 4500 => pixel <= "000000";
      when 4501 => pixel <= "000000";
      when 4502 => pixel <= "000000";
      when 4503 => pixel <= "000000";
      when 4504 => pixel <= "000000";
      when 4505 => pixel <= "000000";
      when 4506 => pixel <= "000000";
      when 4507 => pixel <= "000000";
      when 4508 => pixel <= "000000";
      when 4509 => pixel <= "000000";
      when 4510 => pixel <= "000000";
      when 4511 => pixel <= "000000";
      when 4512 => pixel <= "000000";
      when 4513 => pixel <= "000000";
      when 4514 => pixel <= "000000";
      when 4515 => pixel <= "000000";
      when 4516 => pixel <= "000000";
      when 4517 => pixel <= "000000";
      when 4518 => pixel <= "000000";
      when 4519 => pixel <= "000000";
      when 4520 => pixel <= "000000";
      when 4521 => pixel <= "000000";
      when 4522 => pixel <= "000000";
      when 4523 => pixel <= "000000";
      when 4524 => pixel <= "000000";
      when 4525 => pixel <= "000000";
      when 4526 => pixel <= "000000";
      when 4527 => pixel <= "000000";
      when 4528 => pixel <= "000000";
      when 4529 => pixel <= "000000";
      when 4530 => pixel <= "000000";
      when 4531 => pixel <= "000000";
      when 4532 => pixel <= "000000";
      when 4533 => pixel <= "000000";
      when 4534 => pixel <= "000000";
      when 4535 => pixel <= "000000";
      when 4536 => pixel <= "000000";
      when 4537 => pixel <= "000000";
      when 4538 => pixel <= "000000";
      when 4539 => pixel <= "000000";
      when 4540 => pixel <= "000000";
      when 4541 => pixel <= "000000";
      when 4542 => pixel <= "000000";
      when 4543 => pixel <= "000000";
      when 4544 => pixel <= "000000";
      when 4545 => pixel <= "000000";
      when 4546 => pixel <= "000000";
      when 4547 => pixel <= "000000";
      when 4548 => pixel <= "000000";
      when 4549 => pixel <= "000000";
      when 4550 => pixel <= "000000";
      when 4551 => pixel <= "000000";
      when 4552 => pixel <= "000000";
      when 4553 => pixel <= "000000";
      when 4554 => pixel <= "000000";
      when 4555 => pixel <= "000000";
      when 4556 => pixel <= "000000";
      when 4557 => pixel <= "000000";
      when 4558 => pixel <= "000000";
      when 4559 => pixel <= "000000";
      when 4560 => pixel <= "000000";
      when 4561 => pixel <= "000000";
      when 4562 => pixel <= "000000";
      when 4563 => pixel <= "000000";
      when 4564 => pixel <= "000000";
      when 4565 => pixel <= "000000";
      when 4566 => pixel <= "000000";
      when 4567 => pixel <= "000000";
      when 4568 => pixel <= "000000";
      when 4569 => pixel <= "000000";
      when 4570 => pixel <= "000000";
      when 4571 => pixel <= "000000";
      when 4572 => pixel <= "000000";
      when 4573 => pixel <= "000000";
      when 4574 => pixel <= "000000";
      when 4575 => pixel <= "000000";
      when 4576 => pixel <= "000000";
      when 4577 => pixel <= "000000";
      when 4578 => pixel <= "000000";
      when 4579 => pixel <= "000000";
      when 4580 => pixel <= "000000";
      when 4581 => pixel <= "000000";
      when 4582 => pixel <= "000000";
      when 4583 => pixel <= "000000";
      when 4584 => pixel <= "000000";
      when 4585 => pixel <= "000000";
      when 4586 => pixel <= "000000";
      when 4587 => pixel <= "000000";
      when 4588 => pixel <= "000000";
      when 4589 => pixel <= "000000";
      when 4590 => pixel <= "000000";
      when 4591 => pixel <= "000000";
      when 4592 => pixel <= "000000";
      when 4593 => pixel <= "000000";
      when 4594 => pixel <= "000000";
      when 4595 => pixel <= "000000";
      when 4596 => pixel <= "000000";
      when 4597 => pixel <= "000000";
      when 4598 => pixel <= "000000";
      when 4599 => pixel <= "000000";
      when 4600 => pixel <= "000000";
      when 4601 => pixel <= "000000";
      when 4602 => pixel <= "000000";
      when 4603 => pixel <= "000000";
      when 4604 => pixel <= "000000";
      when 4605 => pixel <= "000000";
      when 4606 => pixel <= "000000";
      when 4607 => pixel <= "000000";
      when 4608 => pixel <= "000000";
      when 4609 => pixel <= "000000";
      when 4610 => pixel <= "000000";
      when 4611 => pixel <= "000000";
      when 4612 => pixel <= "000000";
      when 4613 => pixel <= "000000";
      when 4614 => pixel <= "000000";
      when 4615 => pixel <= "000000";
      when 4616 => pixel <= "000000";
      when 4617 => pixel <= "000000";
      when 4618 => pixel <= "000000";
      when 4619 => pixel <= "000000";
      when 4620 => pixel <= "000000";
      when 4621 => pixel <= "000000";
      when 4622 => pixel <= "000000";
      when 4623 => pixel <= "000000";
      when 4624 => pixel <= "000000";
      when 4625 => pixel <= "000000";
      when 4626 => pixel <= "000000";
      when 4627 => pixel <= "000000";
      when 4628 => pixel <= "000000";
      when 4629 => pixel <= "000000";
      when 4630 => pixel <= "000000";
      when 4631 => pixel <= "000000";
      when 4632 => pixel <= "000000";
      when 4633 => pixel <= "000000";
      when 4634 => pixel <= "000000";
      when 4635 => pixel <= "000000";
      when 4636 => pixel <= "000000";
      when 4637 => pixel <= "000000";
      when 4638 => pixel <= "000000";
      when 4639 => pixel <= "000000";
      when 4640 => pixel <= "000000";
      when 4641 => pixel <= "000000";
      when 4642 => pixel <= "000000";
      when 4643 => pixel <= "000000";
      when 4644 => pixel <= "000000";
      when 4645 => pixel <= "000000";
      when 4646 => pixel <= "000000";
      when 4647 => pixel <= "000000";
      when 4648 => pixel <= "000000";
      when 4649 => pixel <= "000000";
      when 4650 => pixel <= "000000";
      when 4651 => pixel <= "000000";
      when 4652 => pixel <= "000000";
      when 4653 => pixel <= "000000";
      when 4654 => pixel <= "000000";
      when 4655 => pixel <= "000000";
      when 4656 => pixel <= "000000";
      when 4657 => pixel <= "000000";
      when 4658 => pixel <= "000000";
      when 4659 => pixel <= "000000";
      when 4660 => pixel <= "000000";
      when 4661 => pixel <= "000000";
      when 4662 => pixel <= "000000";
      when 4663 => pixel <= "000000";
      when 4664 => pixel <= "000000";
      when 4665 => pixel <= "000000";
      when 4666 => pixel <= "000000";
      when 4667 => pixel <= "000000";
      when 4668 => pixel <= "000000";
      when 4669 => pixel <= "000000";
      when 4670 => pixel <= "000000";
      when 4671 => pixel <= "000000";
      when 4672 => pixel <= "000000";
      when 4673 => pixel <= "000000";
      when 4674 => pixel <= "000000";
      when 4675 => pixel <= "000000";
      when 4676 => pixel <= "000000";
      when 4677 => pixel <= "000000";
      when 4678 => pixel <= "000000";
      when 4679 => pixel <= "000000";
      when 4680 => pixel <= "000000";
      when 4681 => pixel <= "000000";
      when 4682 => pixel <= "000000";
      when 4683 => pixel <= "000000";
      when 4684 => pixel <= "000000";
      when 4685 => pixel <= "000000";
      when 4686 => pixel <= "000000";
      when 4687 => pixel <= "000000";
      when 4688 => pixel <= "000000";
      when 4689 => pixel <= "000000";
      when 4690 => pixel <= "000000";
      when 4691 => pixel <= "000000";
      when 4692 => pixel <= "000000";
      when 4693 => pixel <= "000000";
      when 4694 => pixel <= "000000";
      when 4695 => pixel <= "000000";
      when 4696 => pixel <= "000000";
      when 4697 => pixel <= "000000";
      when 4698 => pixel <= "000000";
      when 4699 => pixel <= "000000";
      when 4700 => pixel <= "000000";
      when 4701 => pixel <= "000000";
      when 4702 => pixel <= "000000";
      when 4703 => pixel <= "000000";
      when 4704 => pixel <= "000000";
      when 4705 => pixel <= "000000";
      when 4706 => pixel <= "000000";
      when 4707 => pixel <= "000000";
      when 4708 => pixel <= "000000";
      when 4709 => pixel <= "000000";
      when 4710 => pixel <= "000000";
      when 4711 => pixel <= "000000";
      when 4712 => pixel <= "000000";
      when 4713 => pixel <= "000000";
      when 4714 => pixel <= "000000";
      when 4715 => pixel <= "000000";
      when 4716 => pixel <= "000000";
      when 4717 => pixel <= "000000";
      when 4718 => pixel <= "000000";
      when 4719 => pixel <= "000000";
      when 4720 => pixel <= "000000";
      when 4721 => pixel <= "000000";
      when 4722 => pixel <= "000000";
      when 4723 => pixel <= "000000";
      when 4724 => pixel <= "000000";
      when 4725 => pixel <= "000000";
      when 4726 => pixel <= "000000";
      when 4727 => pixel <= "000000";
      when 4728 => pixel <= "000000";
      when 4729 => pixel <= "000000";
      when 4730 => pixel <= "000000";
      when 4731 => pixel <= "000000";
      when 4732 => pixel <= "000000";
      when 4733 => pixel <= "000000";
      when 4734 => pixel <= "000000";
      when 4735 => pixel <= "000000";
      when 4736 => pixel <= "000000";
      when 4737 => pixel <= "000000";
      when 4738 => pixel <= "000000";
      when 4739 => pixel <= "000000";
      when 4740 => pixel <= "000000";
      when 4741 => pixel <= "000000";
      when 4742 => pixel <= "000000";
      when 4743 => pixel <= "000000";
      when 4744 => pixel <= "000000";
      when 4745 => pixel <= "000000";
      when 4746 => pixel <= "000000";
      when 4747 => pixel <= "000000";
      when 4748 => pixel <= "000000";
      when 4749 => pixel <= "000000";
      when 4750 => pixel <= "000000";
      when 4751 => pixel <= "000000";
      when 4752 => pixel <= "000000";
      when 4753 => pixel <= "000000";
      when 4754 => pixel <= "000000";
      when 4755 => pixel <= "000000";
      when 4756 => pixel <= "000000";
      when 4757 => pixel <= "000000";
      when 4758 => pixel <= "000000";
      when 4759 => pixel <= "000000";
      when 4760 => pixel <= "000000";
      when 4761 => pixel <= "000000";
      when 4762 => pixel <= "000000";
      when 4763 => pixel <= "000000";
      when 4764 => pixel <= "000000";
      when 4765 => pixel <= "000000";
      when 4766 => pixel <= "000000";
      when 4767 => pixel <= "000000";
      when 4768 => pixel <= "000000";
      when 4769 => pixel <= "000000";
      when 4770 => pixel <= "000000";
      when 4771 => pixel <= "000000";
      when 4772 => pixel <= "000000";
      when 4773 => pixel <= "000000";
      when 4774 => pixel <= "000000";
      when 4775 => pixel <= "000000";
      when 4776 => pixel <= "000000";
      when 4777 => pixel <= "000000";
      when 4778 => pixel <= "000000";
      when 4779 => pixel <= "000000";
      when 4780 => pixel <= "000000";
      when 4781 => pixel <= "000000";
      when 4782 => pixel <= "000000";
      when 4783 => pixel <= "000000";
      when 4784 => pixel <= "000000";
      when 4785 => pixel <= "000000";
      when 4786 => pixel <= "000000";
      when 4787 => pixel <= "000000";
      when 4788 => pixel <= "000000";
      when 4789 => pixel <= "000000";
      when 4790 => pixel <= "000000";
      when 4791 => pixel <= "000000";
      when 4792 => pixel <= "000000";
      when 4793 => pixel <= "000000";
      when 4794 => pixel <= "000000";
      when 4795 => pixel <= "000000";
      when 4796 => pixel <= "000000";
      when 4797 => pixel <= "000000";
      when 4798 => pixel <= "000000";
      when 4799 => pixel <= "000000";
      when 4800 => pixel <= "000000";
      when 4801 => pixel <= "000000";
      when 4802 => pixel <= "000000";
      when 4803 => pixel <= "000000";
      when 4804 => pixel <= "000000";
      when 4805 => pixel <= "000000";
      when 4806 => pixel <= "000000";
      when 4807 => pixel <= "000000";
      when 4808 => pixel <= "000000";
      when 4809 => pixel <= "000000";
      when 4810 => pixel <= "000000";
      when 4811 => pixel <= "000000";
      when 4812 => pixel <= "000000";
      when 4813 => pixel <= "000000";
      when 4814 => pixel <= "000000";
      when 4815 => pixel <= "000000";
      when 4816 => pixel <= "000000";
      when 4817 => pixel <= "000000";
      when 4818 => pixel <= "000000";
      when 4819 => pixel <= "000000";
      when 4820 => pixel <= "000000";
      when 4821 => pixel <= "000000";
      when 4822 => pixel <= "000000";
      when 4823 => pixel <= "000000";
      when 4824 => pixel <= "000000";
      when 4825 => pixel <= "000000";
      when 4826 => pixel <= "000000";
      when 4827 => pixel <= "000000";
      when 4828 => pixel <= "000000";
      when 4829 => pixel <= "000000";
      when 4830 => pixel <= "000000";
      when 4831 => pixel <= "000000";
      when 4832 => pixel <= "000000";
      when 4833 => pixel <= "000000";
      when 4834 => pixel <= "000000";
      when 4835 => pixel <= "000000";
      when 4836 => pixel <= "000000";
      when 4837 => pixel <= "000000";
      when 4838 => pixel <= "000000";
      when 4839 => pixel <= "000000";
      when 4840 => pixel <= "000000";
      when 4841 => pixel <= "000000";
      when 4842 => pixel <= "000000";
      when 4843 => pixel <= "000000";
      when 4844 => pixel <= "000000";
      when 4845 => pixel <= "000000";
      when 4846 => pixel <= "000000";
      when 4847 => pixel <= "000000";
      when 4848 => pixel <= "000000";
      when 4849 => pixel <= "000000";
      when 4850 => pixel <= "000000";
      when 4851 => pixel <= "000000";
      when 4852 => pixel <= "000000";
      when 4853 => pixel <= "000000";
      when 4854 => pixel <= "000000";
      when 4855 => pixel <= "000000";
      when 4856 => pixel <= "000000";
      when 4857 => pixel <= "000000";
      when 4858 => pixel <= "000000";
      when 4859 => pixel <= "000000";
      when 4860 => pixel <= "000000";
      when 4861 => pixel <= "000000";
      when 4862 => pixel <= "000000";
      when 4863 => pixel <= "000000";
      when 4864 => pixel <= "000000";
      when 4865 => pixel <= "000000";
      when 4866 => pixel <= "000000";
      when 4867 => pixel <= "000000";
      when 4868 => pixel <= "000000";
      when 4869 => pixel <= "000000";
      when 4870 => pixel <= "000000";
      when 4871 => pixel <= "000000";
      when 4872 => pixel <= "000000";
      when 4873 => pixel <= "000000";
      when 4874 => pixel <= "000000";
      when 4875 => pixel <= "000000";
      when 4876 => pixel <= "000000";
      when 4877 => pixel <= "000000";
      when 4878 => pixel <= "000000";
      when 4879 => pixel <= "000000";
      when 4880 => pixel <= "000000";
      when 4881 => pixel <= "000000";
      when 4882 => pixel <= "000000";
      when 4883 => pixel <= "000000";
      when 4884 => pixel <= "000000";
      when 4885 => pixel <= "000000";
      when 4886 => pixel <= "000000";
      when 4887 => pixel <= "000000";
      when 4888 => pixel <= "000000";
      when 4889 => pixel <= "000000";
      when 4890 => pixel <= "000000";
      when 4891 => pixel <= "000000";
      when 4892 => pixel <= "000000";
      when 4893 => pixel <= "000000";
      when 4894 => pixel <= "000000";
      when 4895 => pixel <= "000000";
      when 4896 => pixel <= "000000";
      when 4897 => pixel <= "000000";
      when 4898 => pixel <= "000000";
      when 4899 => pixel <= "000000";
      when 4900 => pixel <= "000000";
      when 4901 => pixel <= "000000";
      when 4902 => pixel <= "000000";
      when 4903 => pixel <= "000000";
      when 4904 => pixel <= "000000";
      when 4905 => pixel <= "000000";
      when 4906 => pixel <= "000000";
      when 4907 => pixel <= "000000";
      when 4908 => pixel <= "000000";
      when 4909 => pixel <= "000000";
      when 4910 => pixel <= "000000";
      when 4911 => pixel <= "000000";
      when 4912 => pixel <= "000000";
      when 4913 => pixel <= "000000";
      when 4914 => pixel <= "000000";
      when 4915 => pixel <= "000000";
      when 4916 => pixel <= "000000";
      when 4917 => pixel <= "000000";
      when 4918 => pixel <= "000000";
      when 4919 => pixel <= "000000";
      when 4920 => pixel <= "000000";
      when 4921 => pixel <= "000000";
      when 4922 => pixel <= "000000";
      when 4923 => pixel <= "000000";
      when 4924 => pixel <= "000000";
      when 4925 => pixel <= "000000";
      when 4926 => pixel <= "000000";
      when 4927 => pixel <= "000000";
      when 4928 => pixel <= "000000";
      when 4929 => pixel <= "000000";
      when 4930 => pixel <= "000000";
      when 4931 => pixel <= "000000";
      when 4932 => pixel <= "000000";
      when 4933 => pixel <= "000000";
      when 4934 => pixel <= "000000";
      when 4935 => pixel <= "000000";
      when 4936 => pixel <= "000000";
      when 4937 => pixel <= "000000";
      when 4938 => pixel <= "000000";
      when 4939 => pixel <= "000000";
      when 4940 => pixel <= "000000";
      when 4941 => pixel <= "000000";
      when 4942 => pixel <= "000000";
      when 4943 => pixel <= "000000";
      when 4944 => pixel <= "000000";
      when 4945 => pixel <= "000000";
      when 4946 => pixel <= "000000";
      when 4947 => pixel <= "000000";
      when 4948 => pixel <= "000000";
      when 4949 => pixel <= "000000";
      when 4950 => pixel <= "000000";
      when 4951 => pixel <= "000000";
      when 4952 => pixel <= "000000";
      when 4953 => pixel <= "000000";
      when 4954 => pixel <= "000000";
      when 4955 => pixel <= "000000";
      when 4956 => pixel <= "000000";
      when 4957 => pixel <= "000000";
      when 4958 => pixel <= "000000";
      when 4959 => pixel <= "000000";
      when 4960 => pixel <= "000000";
      when 4961 => pixel <= "000000";
      when 4962 => pixel <= "000000";
      when 4963 => pixel <= "000000";
      when 4964 => pixel <= "000000";
      when 4965 => pixel <= "000000";
      when 4966 => pixel <= "000000";
      when 4967 => pixel <= "000000";
      when 4968 => pixel <= "000000";
      when 4969 => pixel <= "000000";
      when 4970 => pixel <= "000000";
      when 4971 => pixel <= "000000";
      when 4972 => pixel <= "000000";
      when 4973 => pixel <= "000000";
      when 4974 => pixel <= "000000";
      when 4975 => pixel <= "000000";
      when 4976 => pixel <= "000000";
      when 4977 => pixel <= "000000";
      when 4978 => pixel <= "000000";
      when 4979 => pixel <= "000000";
      when 4980 => pixel <= "000000";
      when 4981 => pixel <= "000000";
      when 4982 => pixel <= "000000";
      when 4983 => pixel <= "000000";
      when 4984 => pixel <= "000000";
      when 4985 => pixel <= "000000";
      when 4986 => pixel <= "000000";
      when 4987 => pixel <= "000000";
      when 4988 => pixel <= "000000";
      when 4989 => pixel <= "000000";
      when 4990 => pixel <= "000000";
      when 4991 => pixel <= "000000";
      when 4992 => pixel <= "000000";
      when 4993 => pixel <= "000000";
      when 4994 => pixel <= "000000";
      when 4995 => pixel <= "000000";
      when 4996 => pixel <= "000000";
      when 4997 => pixel <= "000000";
      when 4998 => pixel <= "000000";
      when 4999 => pixel <= "000000";
      when 5000 => pixel <= "000000";
      when 5001 => pixel <= "000000";
      when 5002 => pixel <= "000000";
      when 5003 => pixel <= "000000";
      when 5004 => pixel <= "000000";
      when 5005 => pixel <= "000000";
      when 5006 => pixel <= "000000";
      when 5007 => pixel <= "000000";
      when 5008 => pixel <= "000000";
      when 5009 => pixel <= "000000";
      when 5010 => pixel <= "000000";
      when 5011 => pixel <= "000000";
      when 5012 => pixel <= "000000";
      when 5013 => pixel <= "000000";
      when 5014 => pixel <= "000000";
      when 5015 => pixel <= "000000";
      when 5016 => pixel <= "000000";
      when 5017 => pixel <= "000000";
      when 5018 => pixel <= "000000";
      when 5019 => pixel <= "000000";
      when 5020 => pixel <= "000000";
      when 5021 => pixel <= "000000";
      when 5022 => pixel <= "000000";
      when 5023 => pixel <= "000000";
      when 5024 => pixel <= "000000";
      when 5025 => pixel <= "000000";
      when 5026 => pixel <= "000000";
      when 5027 => pixel <= "000000";
      when 5028 => pixel <= "000000";
      when 5029 => pixel <= "000000";
      when 5030 => pixel <= "000000";
      when 5031 => pixel <= "000000";
      when 5032 => pixel <= "000000";
      when 5033 => pixel <= "000000";
      when 5034 => pixel <= "000000";
      when 5035 => pixel <= "000000";
      when 5036 => pixel <= "000000";
      when 5037 => pixel <= "000000";
      when 5038 => pixel <= "000000";
      when 5039 => pixel <= "000000";
      when 5040 => pixel <= "000000";
      when 5041 => pixel <= "000000";
      when 5042 => pixel <= "000000";
      when 5043 => pixel <= "000000";
      when 5044 => pixel <= "000000";
      when 5045 => pixel <= "000000";
      when 5046 => pixel <= "000000";
      when 5047 => pixel <= "000000";
      when 5048 => pixel <= "000000";
      when 5049 => pixel <= "000000";
      when 5050 => pixel <= "000000";
      when 5051 => pixel <= "000000";
      when 5052 => pixel <= "000000";
      when 5053 => pixel <= "000000";
      when 5054 => pixel <= "000000";
      when 5055 => pixel <= "000000";
      when 5056 => pixel <= "000000";
      when 5057 => pixel <= "000000";
      when 5058 => pixel <= "000000";
      when 5059 => pixel <= "000000";
      when 5060 => pixel <= "000000";
      when 5061 => pixel <= "000000";
      when 5062 => pixel <= "000000";
      when 5063 => pixel <= "000000";
      when 5064 => pixel <= "000000";
      when 5065 => pixel <= "000000";
      when 5066 => pixel <= "000000";
      when 5067 => pixel <= "000000";
      when 5068 => pixel <= "000000";
      when 5069 => pixel <= "000000";
      when 5070 => pixel <= "000000";
      when 5071 => pixel <= "000000";
      when 5072 => pixel <= "000000";
      when 5073 => pixel <= "000000";
      when 5074 => pixel <= "000000";
      when 5075 => pixel <= "000000";
      when 5076 => pixel <= "000000";
      when 5077 => pixel <= "000000";
      when 5078 => pixel <= "000000";
      when 5079 => pixel <= "000000";
      when 5080 => pixel <= "000000";
      when 5081 => pixel <= "000000";
      when 5082 => pixel <= "000000";
      when 5083 => pixel <= "000000";
      when 5084 => pixel <= "000000";
      when 5085 => pixel <= "000000";
      when 5086 => pixel <= "000000";
      when 5087 => pixel <= "000000";
      when 5088 => pixel <= "000000";
      when 5089 => pixel <= "000000";
      when 5090 => pixel <= "000000";
      when 5091 => pixel <= "000000";
      when 5092 => pixel <= "000000";
      when 5093 => pixel <= "000000";
      when 5094 => pixel <= "000000";
      when 5095 => pixel <= "000000";
      when 5096 => pixel <= "000000";
      when 5097 => pixel <= "000000";
      when 5098 => pixel <= "000000";
      when 5099 => pixel <= "000000";
      when 5100 => pixel <= "000000";
      when 5101 => pixel <= "000000";
      when 5102 => pixel <= "000000";
      when 5103 => pixel <= "000000";
      when 5104 => pixel <= "000000";
      when 5105 => pixel <= "000000";
      when 5106 => pixel <= "000000";
      when 5107 => pixel <= "000000";
      when 5108 => pixel <= "000000";
      when 5109 => pixel <= "000000";
      when 5110 => pixel <= "000000";
      when 5111 => pixel <= "000000";
      when 5112 => pixel <= "000000";
      when 5113 => pixel <= "000000";
      when 5114 => pixel <= "000000";
      when 5115 => pixel <= "000000";
      when 5116 => pixel <= "000000";
      when 5117 => pixel <= "000000";
      when 5118 => pixel <= "000000";
      when 5119 => pixel <= "000000";
      when 5120 => pixel <= "000000";
      when 5121 => pixel <= "000000";
      when 5122 => pixel <= "000000";
      when 5123 => pixel <= "000000";
      when 5124 => pixel <= "000000";
      when 5125 => pixel <= "000000";
      when 5126 => pixel <= "000000";
      when 5127 => pixel <= "000000";
      when 5128 => pixel <= "000000";
      when 5129 => pixel <= "000000";
      when 5130 => pixel <= "000000";
      when 5131 => pixel <= "000000";
      when 5132 => pixel <= "000000";
      when 5133 => pixel <= "000000";
      when 5134 => pixel <= "000000";
      when 5135 => pixel <= "000000";
      when 5136 => pixel <= "000000";
      when 5137 => pixel <= "000000";
      when 5138 => pixel <= "000000";
      when 5139 => pixel <= "000000";
      when 5140 => pixel <= "000000";
      when 5141 => pixel <= "000000";
      when 5142 => pixel <= "000000";
      when 5143 => pixel <= "000000";
      when 5144 => pixel <= "000000";
      when 5145 => pixel <= "000000";
      when 5146 => pixel <= "000000";
      when 5147 => pixel <= "000000";
      when 5148 => pixel <= "000000";
      when 5149 => pixel <= "000000";
      when 5150 => pixel <= "000000";
      when 5151 => pixel <= "000000";
      when 5152 => pixel <= "000000";
      when 5153 => pixel <= "000000";
      when 5154 => pixel <= "000000";
      when 5155 => pixel <= "000000";
      when 5156 => pixel <= "000000";
      when 5157 => pixel <= "000000";
      when 5158 => pixel <= "000000";
      when 5159 => pixel <= "000000";
      when 5160 => pixel <= "000000";
      when 5161 => pixel <= "000000";
      when 5162 => pixel <= "000000";
      when 5163 => pixel <= "000000";
      when 5164 => pixel <= "000000";
      when 5165 => pixel <= "000000";
      when 5166 => pixel <= "000000";
      when 5167 => pixel <= "000000";
      when 5168 => pixel <= "000000";
      when 5169 => pixel <= "000000";
      when 5170 => pixel <= "000000";
      when 5171 => pixel <= "000000";
      when 5172 => pixel <= "000000";
      when 5173 => pixel <= "000000";
      when 5174 => pixel <= "000000";
      when 5175 => pixel <= "000000";
      when 5176 => pixel <= "000000";
      when 5177 => pixel <= "000000";
      when 5178 => pixel <= "000000";
      when 5179 => pixel <= "000000";
      when 5180 => pixel <= "000000";
      when 5181 => pixel <= "000000";
      when 5182 => pixel <= "000000";
      when 5183 => pixel <= "000000";
      when 5184 => pixel <= "000000";
      when 5185 => pixel <= "000000";
      when 5186 => pixel <= "000000";
      when 5187 => pixel <= "000000";
      when 5188 => pixel <= "000000";
      when 5189 => pixel <= "000000";
      when 5190 => pixel <= "000000";
      when 5191 => pixel <= "000000";
      when 5192 => pixel <= "000000";
      when 5193 => pixel <= "000000";
      when 5194 => pixel <= "000000";
      when 5195 => pixel <= "000000";
      when 5196 => pixel <= "000000";
      when 5197 => pixel <= "000000";
      when 5198 => pixel <= "000000";
      when 5199 => pixel <= "000000";
      when 5200 => pixel <= "000000";
      when 5201 => pixel <= "000000";
      when 5202 => pixel <= "000000";
      when 5203 => pixel <= "000000";
      when 5204 => pixel <= "000000";
      when 5205 => pixel <= "000000";
      when 5206 => pixel <= "000000";
      when 5207 => pixel <= "000000";
      when 5208 => pixel <= "000000";
      when 5209 => pixel <= "000000";
      when 5210 => pixel <= "000000";
      when 5211 => pixel <= "000000";
      when 5212 => pixel <= "000000";
      when 5213 => pixel <= "000000";
      when 5214 => pixel <= "000000";
      when 5215 => pixel <= "000000";
      when 5216 => pixel <= "000000";
      when 5217 => pixel <= "000000";
      when 5218 => pixel <= "000000";
      when 5219 => pixel <= "000000";
      when 5220 => pixel <= "000000";
      when 5221 => pixel <= "000000";
      when 5222 => pixel <= "000000";
      when 5223 => pixel <= "000000";
      when 5224 => pixel <= "000000";
      when 5225 => pixel <= "000000";
      when 5226 => pixel <= "000000";
      when 5227 => pixel <= "000000";
      when 5228 => pixel <= "000000";
      when 5229 => pixel <= "000000";
      when 5230 => pixel <= "000000";
      when 5231 => pixel <= "000000";
      when 5232 => pixel <= "000000";
      when 5233 => pixel <= "000000";
      when 5234 => pixel <= "000000";
      when 5235 => pixel <= "000000";
      when 5236 => pixel <= "000000";
      when 5237 => pixel <= "000000";
      when 5238 => pixel <= "000000";
      when 5239 => pixel <= "000000";
      when 5240 => pixel <= "000000";
      when 5241 => pixel <= "000000";
      when 5242 => pixel <= "000000";
      when 5243 => pixel <= "000000";
      when 5244 => pixel <= "000000";
      when 5245 => pixel <= "000000";
      when 5246 => pixel <= "000000";
      when 5247 => pixel <= "000000";
      when 5248 => pixel <= "000000";
      when 5249 => pixel <= "000000";
      when 5250 => pixel <= "000000";
      when 5251 => pixel <= "000000";
      when 5252 => pixel <= "000000";
      when 5253 => pixel <= "000000";
      when 5254 => pixel <= "000000";
      when 5255 => pixel <= "000000";
      when 5256 => pixel <= "000000";
      when 5257 => pixel <= "000000";
      when 5258 => pixel <= "000000";
      when 5259 => pixel <= "000000";
      when 5260 => pixel <= "000000";
      when 5261 => pixel <= "000000";
      when 5262 => pixel <= "000000";
      when 5263 => pixel <= "000000";
      when 5264 => pixel <= "000000";
      when 5265 => pixel <= "000000";
      when 5266 => pixel <= "000000";
      when 5267 => pixel <= "000000";
      when 5268 => pixel <= "000000";
      when 5269 => pixel <= "000000";
      when 5270 => pixel <= "000000";
      when 5271 => pixel <= "000000";
      when 5272 => pixel <= "000000";
      when 5273 => pixel <= "000000";
      when 5274 => pixel <= "000000";
      when 5275 => pixel <= "000000";
      when 5276 => pixel <= "000000";
      when 5277 => pixel <= "000000";
      when 5278 => pixel <= "000000";
      when 5279 => pixel <= "000000";
      when 5280 => pixel <= "000000";
      when 5281 => pixel <= "000000";
      when 5282 => pixel <= "000000";
      when 5283 => pixel <= "000000";
      when 5284 => pixel <= "000000";
      when 5285 => pixel <= "000000";
      when 5286 => pixel <= "000000";
      when 5287 => pixel <= "000000";
      when 5288 => pixel <= "000000";
      when 5289 => pixel <= "000000";
      when 5290 => pixel <= "000000";
      when 5291 => pixel <= "000000";
      when 5292 => pixel <= "000000";
      when 5293 => pixel <= "000000";
      when 5294 => pixel <= "000000";
      when 5295 => pixel <= "000000";
      when 5296 => pixel <= "000000";
      when 5297 => pixel <= "000000";
      when 5298 => pixel <= "000000";
      when 5299 => pixel <= "000000";
      when 5300 => pixel <= "000000";
      when 5301 => pixel <= "000000";
      when 5302 => pixel <= "000000";
      when 5303 => pixel <= "000000";
      when 5304 => pixel <= "000000";
      when 5305 => pixel <= "000000";
      when 5306 => pixel <= "000000";
      when 5307 => pixel <= "000000";
      when 5308 => pixel <= "000000";
      when 5309 => pixel <= "000000";
      when 5310 => pixel <= "000000";
      when 5311 => pixel <= "000000";
      when 5312 => pixel <= "000000";
      when 5313 => pixel <= "000000";
      when 5314 => pixel <= "000000";
      when 5315 => pixel <= "000000";
      when 5316 => pixel <= "000000";
      when 5317 => pixel <= "000000";
      when 5318 => pixel <= "000000";
      when 5319 => pixel <= "000000";
      when 5320 => pixel <= "000000";
      when 5321 => pixel <= "000000";
      when 5322 => pixel <= "000000";
      when 5323 => pixel <= "000000";
      when 5324 => pixel <= "000000";
      when 5325 => pixel <= "000000";
      when 5326 => pixel <= "000000";
      when 5327 => pixel <= "000000";
      when 5328 => pixel <= "000000";
      when 5329 => pixel <= "000000";
      when 5330 => pixel <= "000000";
      when 5331 => pixel <= "000000";
      when 5332 => pixel <= "000000";
      when 5333 => pixel <= "000000";
      when 5334 => pixel <= "000000";
      when 5335 => pixel <= "000000";
      when 5336 => pixel <= "000000";
      when 5337 => pixel <= "000000";
      when 5338 => pixel <= "000000";
      when 5339 => pixel <= "000000";
      when 5340 => pixel <= "000000";
      when 5341 => pixel <= "000000";
      when 5342 => pixel <= "000000";
      when 5343 => pixel <= "000000";
      when 5344 => pixel <= "000000";
      when 5345 => pixel <= "000000";
      when 5346 => pixel <= "000000";
      when 5347 => pixel <= "000000";
      when 5348 => pixel <= "000000";
      when 5349 => pixel <= "000000";
      when 5350 => pixel <= "000000";
      when 5351 => pixel <= "000000";
      when 5352 => pixel <= "000000";
      when 5353 => pixel <= "000000";
      when 5354 => pixel <= "000000";
      when 5355 => pixel <= "000000";
      when 5356 => pixel <= "000000";
      when 5357 => pixel <= "000000";
      when 5358 => pixel <= "000000";
      when 5359 => pixel <= "000000";
      when 5360 => pixel <= "000000";
      when 5361 => pixel <= "000000";
      when 5362 => pixel <= "000000";
      when 5363 => pixel <= "000000";
      when 5364 => pixel <= "000000";
      when 5365 => pixel <= "000000";
      when 5366 => pixel <= "000000";
      when 5367 => pixel <= "000000";
      when 5368 => pixel <= "000000";
      when 5369 => pixel <= "000000";
      when 5370 => pixel <= "000000";
      when 5371 => pixel <= "000000";
      when 5372 => pixel <= "000000";
      when 5373 => pixel <= "000000";
      when 5374 => pixel <= "000000";
      when 5375 => pixel <= "000000";
      when 5376 => pixel <= "000000";
      when 5377 => pixel <= "000000";
      when 5378 => pixel <= "000000";
      when 5379 => pixel <= "000000";
      when 5380 => pixel <= "000000";
      when 5381 => pixel <= "000000";
      when 5382 => pixel <= "000000";
      when 5383 => pixel <= "000000";
      when 5384 => pixel <= "000000";
      when 5385 => pixel <= "000000";
      when 5386 => pixel <= "000000";
      when 5387 => pixel <= "000000";
      when 5388 => pixel <= "000000";
      when 5389 => pixel <= "000000";
      when 5390 => pixel <= "000000";
      when 5391 => pixel <= "000000";
      when 5392 => pixel <= "000000";
      when 5393 => pixel <= "000000";
      when 5394 => pixel <= "000000";
      when 5395 => pixel <= "000000";
      when 5396 => pixel <= "000000";
      when 5397 => pixel <= "000000";
      when 5398 => pixel <= "000000";
      when 5399 => pixel <= "000000";
      when 5400 => pixel <= "000000";
      when 5401 => pixel <= "000000";
      when 5402 => pixel <= "000000";
      when 5403 => pixel <= "000000";
      when 5404 => pixel <= "000000";
      when 5405 => pixel <= "000000";
      when 5406 => pixel <= "000000";
      when 5407 => pixel <= "000000";
      when 5408 => pixel <= "000000";
      when 5409 => pixel <= "000000";
      when 5410 => pixel <= "000000";
      when 5411 => pixel <= "000000";
      when 5412 => pixel <= "000000";
      when 5413 => pixel <= "000000";
      when 5414 => pixel <= "000000";
      when 5415 => pixel <= "000000";
      when 5416 => pixel <= "000000";
      when 5417 => pixel <= "000000";
      when 5418 => pixel <= "000000";
      when 5419 => pixel <= "000000";
      when 5420 => pixel <= "000000";
      when 5421 => pixel <= "000000";
      when 5422 => pixel <= "000000";
      when 5423 => pixel <= "000000";
      when 5424 => pixel <= "000000";
      when 5425 => pixel <= "000000";
      when 5426 => pixel <= "000000";
      when 5427 => pixel <= "000000";
      when 5428 => pixel <= "000000";
      when 5429 => pixel <= "000000";
      when 5430 => pixel <= "000000";
      when 5431 => pixel <= "000000";
      when 5432 => pixel <= "000000";
      when 5433 => pixel <= "000000";
      when 5434 => pixel <= "000000";
      when 5435 => pixel <= "000000";
      when 5436 => pixel <= "000000";
      when 5437 => pixel <= "000000";
      when 5438 => pixel <= "000000";
      when 5439 => pixel <= "000000";
      when 5440 => pixel <= "000000";
      when 5441 => pixel <= "000000";
      when 5442 => pixel <= "000000";
      when 5443 => pixel <= "000000";
      when 5444 => pixel <= "000000";
      when 5445 => pixel <= "000000";
      when 5446 => pixel <= "000000";
      when 5447 => pixel <= "000000";
      when 5448 => pixel <= "000000";
      when 5449 => pixel <= "000000";
      when 5450 => pixel <= "000000";
      when 5451 => pixel <= "000000";
      when 5452 => pixel <= "000000";
      when 5453 => pixel <= "000000";
      when 5454 => pixel <= "000000";
      when 5455 => pixel <= "000000";
      when 5456 => pixel <= "000000";
      when 5457 => pixel <= "000000";
      when 5458 => pixel <= "000000";
      when 5459 => pixel <= "000000";
      when 5460 => pixel <= "000000";
      when 5461 => pixel <= "000000";
      when 5462 => pixel <= "000000";
      when 5463 => pixel <= "000000";
      when 5464 => pixel <= "000000";
      when 5465 => pixel <= "000000";
      when 5466 => pixel <= "000000";
      when 5467 => pixel <= "000000";
      when 5468 => pixel <= "000000";
      when 5469 => pixel <= "000000";
      when 5470 => pixel <= "000000";
      when 5471 => pixel <= "000000";
      when 5472 => pixel <= "000000";
      when 5473 => pixel <= "000000";
      when 5474 => pixel <= "000000";
      when 5475 => pixel <= "000000";
      when 5476 => pixel <= "000000";
      when 5477 => pixel <= "000000";
      when 5478 => pixel <= "000000";
      when 5479 => pixel <= "000000";
      when 5480 => pixel <= "000000";
      when 5481 => pixel <= "000000";
      when 5482 => pixel <= "000000";
      when 5483 => pixel <= "000000";
      when 5484 => pixel <= "000000";
      when 5485 => pixel <= "000000";
      when 5486 => pixel <= "000000";
      when 5487 => pixel <= "000000";
      when 5488 => pixel <= "000000";
      when 5489 => pixel <= "000000";
      when 5490 => pixel <= "000000";
      when 5491 => pixel <= "000000";
      when 5492 => pixel <= "000000";
      when 5493 => pixel <= "000000";
      when 5494 => pixel <= "000000";
      when 5495 => pixel <= "000000";
      when 5496 => pixel <= "000000";
      when 5497 => pixel <= "000000";
      when 5498 => pixel <= "000000";
      when 5499 => pixel <= "000000";
      when 5500 => pixel <= "000000";
      when 5501 => pixel <= "000000";
      when 5502 => pixel <= "000000";
      when 5503 => pixel <= "000000";
      when 5504 => pixel <= "000000";
      when 5505 => pixel <= "000000";
      when 5506 => pixel <= "000000";
      when 5507 => pixel <= "000000";
      when 5508 => pixel <= "000000";
      when 5509 => pixel <= "000000";
      when 5510 => pixel <= "000000";
      when 5511 => pixel <= "000000";
      when 5512 => pixel <= "000000";
      when 5513 => pixel <= "000000";
      when 5514 => pixel <= "000000";
      when 5515 => pixel <= "000000";
      when 5516 => pixel <= "000000";
      when 5517 => pixel <= "000000";
      when 5518 => pixel <= "000000";
      when 5519 => pixel <= "000000";
      when 5520 => pixel <= "000000";
      when 5521 => pixel <= "000000";
      when 5522 => pixel <= "000000";
      when 5523 => pixel <= "000000";
      when 5524 => pixel <= "000000";
      when 5525 => pixel <= "000000";
      when 5526 => pixel <= "000000";
      when 5527 => pixel <= "000000";
      when 5528 => pixel <= "000000";
      when 5529 => pixel <= "000000";
      when 5530 => pixel <= "000000";
      when 5531 => pixel <= "000000";
      when 5532 => pixel <= "000000";
      when 5533 => pixel <= "000000";
      when 5534 => pixel <= "000000";
      when 5535 => pixel <= "000000";
      when 5536 => pixel <= "000000";
      when 5537 => pixel <= "000000";
      when 5538 => pixel <= "000000";
      when 5539 => pixel <= "000000";
      when 5540 => pixel <= "000000";
      when 5541 => pixel <= "000000";
      when 5542 => pixel <= "000000";
      when 5543 => pixel <= "000000";
      when 5544 => pixel <= "000000";
      when 5545 => pixel <= "000000";
      when 5546 => pixel <= "000000";
      when 5547 => pixel <= "000000";
      when 5548 => pixel <= "000000";
      when 5549 => pixel <= "000000";
      when 5550 => pixel <= "000000";
      when 5551 => pixel <= "000000";
      when 5552 => pixel <= "000000";
      when 5553 => pixel <= "000000";
      when 5554 => pixel <= "000000";
      when 5555 => pixel <= "000000";
      when 5556 => pixel <= "000000";
      when 5557 => pixel <= "000000";
      when 5558 => pixel <= "000000";
      when 5559 => pixel <= "000000";
      when 5560 => pixel <= "000000";
      when 5561 => pixel <= "000000";
      when 5562 => pixel <= "000000";
      when 5563 => pixel <= "000000";
      when 5564 => pixel <= "000000";
      when 5565 => pixel <= "000000";
      when 5566 => pixel <= "000000";
      when 5567 => pixel <= "000000";
      when 5568 => pixel <= "000000";
      when 5569 => pixel <= "000000";
      when 5570 => pixel <= "000000";
      when 5571 => pixel <= "000000";
      when 5572 => pixel <= "000000";
      when 5573 => pixel <= "000000";
      when 5574 => pixel <= "000000";
      when 5575 => pixel <= "000000";
      when 5576 => pixel <= "000000";
      when 5577 => pixel <= "000000";
      when 5578 => pixel <= "000000";
      when 5579 => pixel <= "000000";
      when 5580 => pixel <= "000000";
      when 5581 => pixel <= "000000";
      when 5582 => pixel <= "000000";
      when 5583 => pixel <= "000000";
      when 5584 => pixel <= "000000";
      when 5585 => pixel <= "000000";
      when 5586 => pixel <= "000000";
      when 5587 => pixel <= "000000";
      when 5588 => pixel <= "000000";
      when 5589 => pixel <= "000000";
      when 5590 => pixel <= "000000";
      when 5591 => pixel <= "000000";
      when 5592 => pixel <= "000000";
      when 5593 => pixel <= "000000";
      when 5594 => pixel <= "000000";
      when 5595 => pixel <= "000000";
      when 5596 => pixel <= "000000";
      when 5597 => pixel <= "000000";
      when 5598 => pixel <= "000000";
      when 5599 => pixel <= "000000";
      when 5600 => pixel <= "000000";
      when 5601 => pixel <= "000000";
      when 5602 => pixel <= "000000";
      when 5603 => pixel <= "000000";
      when 5604 => pixel <= "000000";
      when 5605 => pixel <= "000000";
      when 5606 => pixel <= "000000";
      when 5607 => pixel <= "000000";
      when 5608 => pixel <= "000000";
      when 5609 => pixel <= "000000";
      when 5610 => pixel <= "000000";
      when 5611 => pixel <= "000000";
      when 5612 => pixel <= "000000";
      when 5613 => pixel <= "000000";
      when 5614 => pixel <= "000000";
      when 5615 => pixel <= "000000";
      when 5616 => pixel <= "000000";
      when 5617 => pixel <= "000000";
      when 5618 => pixel <= "000000";
      when 5619 => pixel <= "000000";
      when 5620 => pixel <= "000000";
      when 5621 => pixel <= "000000";
      when 5622 => pixel <= "000000";
      when 5623 => pixel <= "000000";
      when 5624 => pixel <= "000000";
      when 5625 => pixel <= "000000";
      when 5626 => pixel <= "000000";
      when 5627 => pixel <= "000000";
      when 5628 => pixel <= "000000";
      when 5629 => pixel <= "000000";
      when 5630 => pixel <= "000000";
      when 5631 => pixel <= "000000";
      when 5632 => pixel <= "000000";
      when 5633 => pixel <= "000000";
      when 5634 => pixel <= "000000";
      when 5635 => pixel <= "000000";
      when 5636 => pixel <= "000000";
      when 5637 => pixel <= "000000";
      when 5638 => pixel <= "000000";
      when 5639 => pixel <= "000000";
      when 5640 => pixel <= "000000";
      when 5641 => pixel <= "000000";
      when 5642 => pixel <= "000000";
      when 5643 => pixel <= "000000";
      when 5644 => pixel <= "000000";
      when 5645 => pixel <= "000000";
      when 5646 => pixel <= "000000";
      when 5647 => pixel <= "000000";
      when 5648 => pixel <= "000000";
      when 5649 => pixel <= "000000";
      when 5650 => pixel <= "000000";
      when 5651 => pixel <= "000000";
      when 5652 => pixel <= "000000";
      when 5653 => pixel <= "000000";
      when 5654 => pixel <= "000000";
      when 5655 => pixel <= "000000";
      when 5656 => pixel <= "000000";
      when 5657 => pixel <= "000000";
      when 5658 => pixel <= "000000";
      when 5659 => pixel <= "000000";
      when 5660 => pixel <= "000000";
      when 5661 => pixel <= "000000";
      when 5662 => pixel <= "000000";
      when 5663 => pixel <= "000000";
      when 5664 => pixel <= "000000";
      when 5665 => pixel <= "000000";
      when 5666 => pixel <= "000000";
      when 5667 => pixel <= "000000";
      when 5668 => pixel <= "000000";
      when 5669 => pixel <= "000000";
      when 5670 => pixel <= "000000";
      when 5671 => pixel <= "000000";
      when 5672 => pixel <= "000000";
      when 5673 => pixel <= "000000";
      when 5674 => pixel <= "000000";
      when 5675 => pixel <= "000000";
      when 5676 => pixel <= "000000";
      when 5677 => pixel <= "000000";
      when 5678 => pixel <= "000000";
      when 5679 => pixel <= "000000";
      when 5680 => pixel <= "000000";
      when 5681 => pixel <= "000000";
      when 5682 => pixel <= "000000";
      when 5683 => pixel <= "000000";
      when 5684 => pixel <= "000000";
      when 5685 => pixel <= "000000";
      when 5686 => pixel <= "000000";
      when 5687 => pixel <= "000000";
      when 5688 => pixel <= "000000";
      when 5689 => pixel <= "000000";
      when 5690 => pixel <= "000000";
      when 5691 => pixel <= "000000";
      when 5692 => pixel <= "000000";
      when 5693 => pixel <= "000000";
      when 5694 => pixel <= "000000";
      when 5695 => pixel <= "000000";
      when 5696 => pixel <= "000000";
      when 5697 => pixel <= "000000";
      when 5698 => pixel <= "000000";
      when 5699 => pixel <= "000000";
      when 5700 => pixel <= "000000";
      when 5701 => pixel <= "000000";
      when 5702 => pixel <= "000000";
      when 5703 => pixel <= "000000";
      when 5704 => pixel <= "000000";
      when 5705 => pixel <= "000000";
      when 5706 => pixel <= "000000";
      when 5707 => pixel <= "000000";
      when 5708 => pixel <= "000000";
      when 5709 => pixel <= "000000";
      when 5710 => pixel <= "000000";
      when 5711 => pixel <= "000000";
      when 5712 => pixel <= "000000";
      when 5713 => pixel <= "000000";
      when 5714 => pixel <= "000000";
      when 5715 => pixel <= "000000";
      when 5716 => pixel <= "000000";
      when 5717 => pixel <= "000000";
      when 5718 => pixel <= "000000";
      when 5719 => pixel <= "000000";
      when 5720 => pixel <= "000000";
      when 5721 => pixel <= "000000";
      when 5722 => pixel <= "000000";
      when 5723 => pixel <= "000000";
      when 5724 => pixel <= "000000";
      when 5725 => pixel <= "000000";
      when 5726 => pixel <= "000000";
      when 5727 => pixel <= "000000";
      when 5728 => pixel <= "000000";
      when 5729 => pixel <= "000000";
      when 5730 => pixel <= "000000";
      when 5731 => pixel <= "000000";
      when 5732 => pixel <= "000000";
      when 5733 => pixel <= "000000";
      when 5734 => pixel <= "000000";
      when 5735 => pixel <= "000000";
      when 5736 => pixel <= "000000";
      when 5737 => pixel <= "000000";
      when 5738 => pixel <= "000000";
      when 5739 => pixel <= "000000";
      when 5740 => pixel <= "000000";
      when 5741 => pixel <= "000000";
      when 5742 => pixel <= "000000";
      when 5743 => pixel <= "000000";
      when 5744 => pixel <= "000000";
      when 5745 => pixel <= "000000";
      when 5746 => pixel <= "000000";
      when 5747 => pixel <= "000000";
      when 5748 => pixel <= "000000";
      when 5749 => pixel <= "000000";
      when 5750 => pixel <= "000000";
      when 5751 => pixel <= "000000";
      when 5752 => pixel <= "000000";
      when 5753 => pixel <= "000000";
      when 5754 => pixel <= "000000";
      when 5755 => pixel <= "000000";
      when 5756 => pixel <= "000000";
      when 5757 => pixel <= "000000";
      when 5758 => pixel <= "000000";
      when 5759 => pixel <= "000000";
      when 5760 => pixel <= "000000";
      when 5761 => pixel <= "000000";
      when 5762 => pixel <= "000000";
      when 5763 => pixel <= "000000";
      when 5764 => pixel <= "000000";
      when 5765 => pixel <= "000000";
      when 5766 => pixel <= "000000";
      when 5767 => pixel <= "000000";
      when 5768 => pixel <= "000000";
      when 5769 => pixel <= "000000";
      when 5770 => pixel <= "000000";
      when 5771 => pixel <= "000000";
      when 5772 => pixel <= "000000";
      when 5773 => pixel <= "000000";
      when 5774 => pixel <= "000000";
      when 5775 => pixel <= "000000";
      when 5776 => pixel <= "000000";
      when 5777 => pixel <= "000000";
      when 5778 => pixel <= "000000";
      when 5779 => pixel <= "000000";
      when 5780 => pixel <= "000000";
      when 5781 => pixel <= "000000";
      when 5782 => pixel <= "000000";
      when 5783 => pixel <= "000000";
      when 5784 => pixel <= "000000";
      when 5785 => pixel <= "000000";
      when 5786 => pixel <= "000000";
      when 5787 => pixel <= "000000";
      when 5788 => pixel <= "000000";
      when 5789 => pixel <= "000000";
      when 5790 => pixel <= "000000";
      when 5791 => pixel <= "000000";
      when 5792 => pixel <= "000000";
      when 5793 => pixel <= "000000";
      when 5794 => pixel <= "000000";
      when 5795 => pixel <= "000000";
      when 5796 => pixel <= "000000";
      when 5797 => pixel <= "000000";
      when 5798 => pixel <= "000000";
      when 5799 => pixel <= "000000";
      when 5800 => pixel <= "000000";
      when 5801 => pixel <= "000000";
      when 5802 => pixel <= "000000";
      when 5803 => pixel <= "000000";
      when 5804 => pixel <= "000000";
      when 5805 => pixel <= "000000";
      when 5806 => pixel <= "000000";
      when 5807 => pixel <= "000000";
      when 5808 => pixel <= "000000";
      when 5809 => pixel <= "000000";
      when 5810 => pixel <= "000000";
      when 5811 => pixel <= "000000";
      when 5812 => pixel <= "000000";
      when 5813 => pixel <= "000000";
      when 5814 => pixel <= "000000";
      when 5815 => pixel <= "000000";
      when 5816 => pixel <= "000000";
      when 5817 => pixel <= "000000";
      when 5818 => pixel <= "000000";
      when 5819 => pixel <= "000000";
      when 5820 => pixel <= "000000";
      when 5821 => pixel <= "000000";
      when 5822 => pixel <= "000000";
      when 5823 => pixel <= "000000";
      when 5824 => pixel <= "000000";
      when 5825 => pixel <= "000000";
      when 5826 => pixel <= "000000";
      when 5827 => pixel <= "000000";
      when 5828 => pixel <= "000000";
      when 5829 => pixel <= "000000";
      when 5830 => pixel <= "000000";
      when 5831 => pixel <= "000000";
      when 5832 => pixel <= "000000";
      when 5833 => pixel <= "000000";
      when 5834 => pixel <= "000000";
      when 5835 => pixel <= "000000";
      when 5836 => pixel <= "000000";
      when 5837 => pixel <= "000000";
      when 5838 => pixel <= "000000";
      when 5839 => pixel <= "000000";
      when 5840 => pixel <= "000000";
      when 5841 => pixel <= "000000";
      when 5842 => pixel <= "000000";
      when 5843 => pixel <= "000000";
      when 5844 => pixel <= "000000";
      when 5845 => pixel <= "000000";
      when 5846 => pixel <= "000000";
      when 5847 => pixel <= "000000";
      when 5848 => pixel <= "000000";
      when 5849 => pixel <= "000000";
      when 5850 => pixel <= "000000";
      when 5851 => pixel <= "000000";
      when 5852 => pixel <= "000000";
      when 5853 => pixel <= "000000";
      when 5854 => pixel <= "000000";
      when 5855 => pixel <= "000000";
      when 5856 => pixel <= "000000";
      when 5857 => pixel <= "000000";
      when 5858 => pixel <= "000000";
      when 5859 => pixel <= "000000";
      when 5860 => pixel <= "000000";
      when 5861 => pixel <= "000000";
      when 5862 => pixel <= "000000";
      when 5863 => pixel <= "000000";
      when 5864 => pixel <= "000000";
      when 5865 => pixel <= "000000";
      when 5866 => pixel <= "000000";
      when 5867 => pixel <= "000000";
      when 5868 => pixel <= "000000";
      when 5869 => pixel <= "000000";
      when 5870 => pixel <= "000000";
      when 5871 => pixel <= "000000";
      when 5872 => pixel <= "000000";
      when 5873 => pixel <= "000000";
      when 5874 => pixel <= "000000";
      when 5875 => pixel <= "000000";
      when 5876 => pixel <= "000000";
      when 5877 => pixel <= "000000";
      when 5878 => pixel <= "000000";
      when 5879 => pixel <= "000000";
      when 5880 => pixel <= "000000";
      when 5881 => pixel <= "000000";
      when 5882 => pixel <= "000000";
      when 5883 => pixel <= "000000";
      when 5884 => pixel <= "000000";
      when 5885 => pixel <= "000000";
      when 5886 => pixel <= "000000";
      when 5887 => pixel <= "000000";
      when 5888 => pixel <= "000000";
      when 5889 => pixel <= "000000";
      when 5890 => pixel <= "000000";
      when 5891 => pixel <= "000000";
      when 5892 => pixel <= "000000";
      when 5893 => pixel <= "000000";
      when 5894 => pixel <= "000000";
      when 5895 => pixel <= "000000";
      when 5896 => pixel <= "000000";
      when 5897 => pixel <= "000000";
      when 5898 => pixel <= "000000";
      when 5899 => pixel <= "000000";
      when 5900 => pixel <= "000000";
      when 5901 => pixel <= "000000";
      when 5902 => pixel <= "000000";
      when 5903 => pixel <= "000000";
      when 5904 => pixel <= "000000";
      when 5905 => pixel <= "000000";
      when 5906 => pixel <= "000000";
      when 5907 => pixel <= "000000";
      when 5908 => pixel <= "000000";
      when 5909 => pixel <= "000000";
      when 5910 => pixel <= "000000";
      when 5911 => pixel <= "000000";
      when 5912 => pixel <= "000000";
      when 5913 => pixel <= "000000";
      when 5914 => pixel <= "000000";
      when 5915 => pixel <= "000000";
      when 5916 => pixel <= "000000";
      when 5917 => pixel <= "000000";
      when 5918 => pixel <= "000000";
      when 5919 => pixel <= "000000";
      when 5920 => pixel <= "000000";
      when 5921 => pixel <= "000000";
      when 5922 => pixel <= "000000";
      when 5923 => pixel <= "000000";
      when 5924 => pixel <= "000000";
      when 5925 => pixel <= "000000";
      when 5926 => pixel <= "000000";
      when 5927 => pixel <= "000000";
      when 5928 => pixel <= "000000";
      when 5929 => pixel <= "000000";
      when 5930 => pixel <= "000000";
      when 5931 => pixel <= "000000";
      when 5932 => pixel <= "000000";
      when 5933 => pixel <= "000000";
      when 5934 => pixel <= "000000";
      when 5935 => pixel <= "000000";
      when 5936 => pixel <= "000000";
      when 5937 => pixel <= "000000";
      when 5938 => pixel <= "000000";
      when 5939 => pixel <= "000000";
      when 5940 => pixel <= "000000";
      when 5941 => pixel <= "000000";
      when 5942 => pixel <= "000000";
      when 5943 => pixel <= "000000";
      when 5944 => pixel <= "000000";
      when 5945 => pixel <= "000000";
      when 5946 => pixel <= "000000";
      when 5947 => pixel <= "000000";
      when 5948 => pixel <= "000000";
      when 5949 => pixel <= "000000";
      when 5950 => pixel <= "000000";
      when 5951 => pixel <= "000000";
      when 5952 => pixel <= "000000";
      when 5953 => pixel <= "000000";
      when 5954 => pixel <= "000000";
      when 5955 => pixel <= "000000";
      when 5956 => pixel <= "000000";
      when 5957 => pixel <= "000000";
      when 5958 => pixel <= "000000";
      when 5959 => pixel <= "000000";
      when 5960 => pixel <= "000000";
      when 5961 => pixel <= "000000";
      when 5962 => pixel <= "000000";
      when 5963 => pixel <= "000000";
      when 5964 => pixel <= "000000";
      when 5965 => pixel <= "000000";
      when 5966 => pixel <= "000000";
      when 5967 => pixel <= "000000";
      when 5968 => pixel <= "000000";
      when 5969 => pixel <= "000000";
      when 5970 => pixel <= "000000";
      when 5971 => pixel <= "000000";
      when 5972 => pixel <= "000000";
      when 5973 => pixel <= "000000";
      when 5974 => pixel <= "000000";
      when 5975 => pixel <= "000000";
      when 5976 => pixel <= "000000";
      when 5977 => pixel <= "000000";
      when 5978 => pixel <= "000000";
      when 5979 => pixel <= "000000";
      when 5980 => pixel <= "000000";
      when 5981 => pixel <= "000000";
      when 5982 => pixel <= "000000";
      when 5983 => pixel <= "000000";
      when 5984 => pixel <= "000000";
      when 5985 => pixel <= "000000";
      when 5986 => pixel <= "000000";
      when 5987 => pixel <= "000000";
      when 5988 => pixel <= "000000";
      when 5989 => pixel <= "000000";
      when 5990 => pixel <= "000000";
      when 5991 => pixel <= "000000";
      when 5992 => pixel <= "000000";
      when 5993 => pixel <= "000000";
      when 5994 => pixel <= "000000";
      when 5995 => pixel <= "000000";
      when 5996 => pixel <= "000000";
      when 5997 => pixel <= "000000";
      when 5998 => pixel <= "000000";
      when 5999 => pixel <= "000000";
      when 6000 => pixel <= "000000";
      when 6001 => pixel <= "000000";
      when 6002 => pixel <= "000000";
      when 6003 => pixel <= "000000";
      when 6004 => pixel <= "000000";
      when 6005 => pixel <= "000000";
      when 6006 => pixel <= "000000";
      when 6007 => pixel <= "000000";
      when 6008 => pixel <= "000000";
      when 6009 => pixel <= "000000";
      when 6010 => pixel <= "000000";
      when 6011 => pixel <= "000000";
      when 6012 => pixel <= "000000";
      when 6013 => pixel <= "000000";
      when 6014 => pixel <= "000000";
      when 6015 => pixel <= "000000";
      when 6016 => pixel <= "000000";
      when 6017 => pixel <= "000000";
      when 6018 => pixel <= "000000";
      when 6019 => pixel <= "000000";
      when 6020 => pixel <= "000000";
      when 6021 => pixel <= "000000";
      when 6022 => pixel <= "000000";
      when 6023 => pixel <= "000000";
      when 6024 => pixel <= "000000";
      when 6025 => pixel <= "000000";
      when 6026 => pixel <= "000000";
      when 6027 => pixel <= "000000";
      when 6028 => pixel <= "000000";
      when 6029 => pixel <= "000000";
      when 6030 => pixel <= "000000";
      when 6031 => pixel <= "000000";
      when 6032 => pixel <= "000000";
      when 6033 => pixel <= "000000";
      when 6034 => pixel <= "000000";
      when 6035 => pixel <= "000000";
      when 6036 => pixel <= "000000";
      when 6037 => pixel <= "000000";
      when 6038 => pixel <= "000000";
      when 6039 => pixel <= "000000";
      when 6040 => pixel <= "000000";
      when 6041 => pixel <= "000000";
      when 6042 => pixel <= "000000";
      when 6043 => pixel <= "000000";
      when 6044 => pixel <= "000000";
      when 6045 => pixel <= "000000";
      when 6046 => pixel <= "000000";
      when 6047 => pixel <= "000000";
      when 6048 => pixel <= "000000";
      when 6049 => pixel <= "000000";
      when 6050 => pixel <= "000000";
      when 6051 => pixel <= "000000";
      when 6052 => pixel <= "000000";
      when 6053 => pixel <= "000000";
      when 6054 => pixel <= "000000";
      when 6055 => pixel <= "000000";
      when 6056 => pixel <= "000000";
      when 6057 => pixel <= "000000";
      when 6058 => pixel <= "000000";
      when 6059 => pixel <= "000000";
      when 6060 => pixel <= "000000";
      when 6061 => pixel <= "000000";
      when 6062 => pixel <= "000000";
      when 6063 => pixel <= "000000";
      when 6064 => pixel <= "000000";
      when 6065 => pixel <= "000000";
      when 6066 => pixel <= "000000";
      when 6067 => pixel <= "000000";
      when 6068 => pixel <= "000000";
      when 6069 => pixel <= "000000";
      when 6070 => pixel <= "000000";
      when 6071 => pixel <= "000000";
      when 6072 => pixel <= "000000";
      when 6073 => pixel <= "000000";
      when 6074 => pixel <= "000000";
      when 6075 => pixel <= "000000";
      when 6076 => pixel <= "000000";
      when 6077 => pixel <= "000000";
      when 6078 => pixel <= "000000";
      when 6079 => pixel <= "000000";
      when 6080 => pixel <= "000000";
      when 6081 => pixel <= "000000";
      when 6082 => pixel <= "000000";
      when 6083 => pixel <= "000000";
      when 6084 => pixel <= "000000";
      when 6085 => pixel <= "000000";
      when 6086 => pixel <= "000000";
      when 6087 => pixel <= "000000";
      when 6088 => pixel <= "000000";
      when 6089 => pixel <= "000000";
      when 6090 => pixel <= "000000";
      when 6091 => pixel <= "000000";
      when 6092 => pixel <= "000000";
      when 6093 => pixel <= "000000";
      when 6094 => pixel <= "000000";
      when 6095 => pixel <= "000000";
      when 6096 => pixel <= "000000";
      when 6097 => pixel <= "000000";
      when 6098 => pixel <= "000000";
      when 6099 => pixel <= "000000";
      when 6100 => pixel <= "000000";
      when 6101 => pixel <= "000000";
      when 6102 => pixel <= "000000";
      when 6103 => pixel <= "000000";
      when 6104 => pixel <= "000000";
      when 6105 => pixel <= "000000";
      when 6106 => pixel <= "000000";
      when 6107 => pixel <= "000000";
      when 6108 => pixel <= "000000";
      when 6109 => pixel <= "000000";
      when 6110 => pixel <= "000000";
      when 6111 => pixel <= "000000";
      when 6112 => pixel <= "000000";
      when 6113 => pixel <= "000000";
      when 6114 => pixel <= "000000";
      when 6115 => pixel <= "000000";
      when 6116 => pixel <= "000000";
      when 6117 => pixel <= "000000";
      when 6118 => pixel <= "000000";
      when 6119 => pixel <= "000000";
      when 6120 => pixel <= "000000";
      when 6121 => pixel <= "000000";
      when 6122 => pixel <= "000000";
      when 6123 => pixel <= "000000";
      when 6124 => pixel <= "000000";
      when 6125 => pixel <= "000000";
      when 6126 => pixel <= "000000";
      when 6127 => pixel <= "000000";
      when 6128 => pixel <= "000000";
      when 6129 => pixel <= "000000";
      when 6130 => pixel <= "000000";
      when 6131 => pixel <= "000000";
      when 6132 => pixel <= "000000";
      when 6133 => pixel <= "000000";
      when 6134 => pixel <= "000000";
      when 6135 => pixel <= "000000";
      when 6136 => pixel <= "000000";
      when 6137 => pixel <= "000000";
      when 6138 => pixel <= "000000";
      when 6139 => pixel <= "000000";
      when 6140 => pixel <= "000000";
      when 6141 => pixel <= "000000";
      when 6142 => pixel <= "000000";
      when 6143 => pixel <= "000000";
      when 6144 => pixel <= "000000";
      when 6145 => pixel <= "000000";
      when 6146 => pixel <= "000000";
      when 6147 => pixel <= "000000";
      when 6148 => pixel <= "000000";
      when 6149 => pixel <= "000000";
      when 6150 => pixel <= "000000";
      when 6151 => pixel <= "000000";
      when 6152 => pixel <= "000000";
      when 6153 => pixel <= "000000";
      when 6154 => pixel <= "000000";
      when 6155 => pixel <= "000000";
      when 6156 => pixel <= "000000";
      when 6157 => pixel <= "000000";
      when 6158 => pixel <= "000000";
      when 6159 => pixel <= "000000";
      when 6160 => pixel <= "000000";
      when 6161 => pixel <= "000000";
      when 6162 => pixel <= "000000";
      when 6163 => pixel <= "000000";
      when 6164 => pixel <= "000000";
      when 6165 => pixel <= "000000";
      when 6166 => pixel <= "000000";
      when 6167 => pixel <= "000000";
      when 6168 => pixel <= "000000";
      when 6169 => pixel <= "000000";
      when 6170 => pixel <= "000000";
      when 6171 => pixel <= "000000";
      when 6172 => pixel <= "000000";
      when 6173 => pixel <= "000000";
      when 6174 => pixel <= "000000";
      when 6175 => pixel <= "000000";
      when 6176 => pixel <= "000000";
      when 6177 => pixel <= "000000";
      when 6178 => pixel <= "000000";
      when 6179 => pixel <= "000000";
      when 6180 => pixel <= "000000";
      when 6181 => pixel <= "000000";
      when 6182 => pixel <= "000000";
      when 6183 => pixel <= "000000";
      when 6184 => pixel <= "000000";
      when 6185 => pixel <= "000000";
      when 6186 => pixel <= "000000";
      when 6187 => pixel <= "000000";
      when 6188 => pixel <= "000000";
      when 6189 => pixel <= "000000";
      when 6190 => pixel <= "000000";
      when 6191 => pixel <= "000000";
      when 6192 => pixel <= "000000";
      when 6193 => pixel <= "000000";
      when 6194 => pixel <= "000000";
      when 6195 => pixel <= "000000";
      when 6196 => pixel <= "000000";
      when 6197 => pixel <= "000000";
      when 6198 => pixel <= "000000";
      when 6199 => pixel <= "000000";
      when 6200 => pixel <= "000000";
      when 6201 => pixel <= "000000";
      when 6202 => pixel <= "000000";
      when 6203 => pixel <= "000000";
      when 6204 => pixel <= "000000";
      when 6205 => pixel <= "000000";
      when 6206 => pixel <= "000000";
      when 6207 => pixel <= "000000";
      when 6208 => pixel <= "000000";
      when 6209 => pixel <= "000000";
      when 6210 => pixel <= "000000";
      when 6211 => pixel <= "000000";
      when 6212 => pixel <= "000000";
      when 6213 => pixel <= "000000";
      when 6214 => pixel <= "000000";
      when 6215 => pixel <= "000000";
      when 6216 => pixel <= "000000";
      when 6217 => pixel <= "000000";
      when 6218 => pixel <= "000000";
      when 6219 => pixel <= "000000";
      when 6220 => pixel <= "000000";
      when 6221 => pixel <= "000000";
      when 6222 => pixel <= "000000";
      when 6223 => pixel <= "000000";
      when 6224 => pixel <= "000000";
      when 6225 => pixel <= "000000";
      when 6226 => pixel <= "000000";
      when 6227 => pixel <= "000000";
      when 6228 => pixel <= "000000";
      when 6229 => pixel <= "000000";
      when 6230 => pixel <= "000000";
      when 6231 => pixel <= "000000";
      when 6232 => pixel <= "000000";
      when 6233 => pixel <= "000000";
      when 6234 => pixel <= "000000";
      when 6235 => pixel <= "000000";
      when 6236 => pixel <= "000000";
      when 6237 => pixel <= "000000";
      when 6238 => pixel <= "000000";
      when 6239 => pixel <= "000000";
      when 6240 => pixel <= "000000";
      when 6241 => pixel <= "000000";
      when 6242 => pixel <= "000000";
      when 6243 => pixel <= "000000";
      when 6244 => pixel <= "000000";
      when 6245 => pixel <= "000000";
      when 6246 => pixel <= "000000";
      when 6247 => pixel <= "000000";
      when 6248 => pixel <= "000000";
      when 6249 => pixel <= "000000";
      when 6250 => pixel <= "000000";
      when 6251 => pixel <= "000000";
      when 6252 => pixel <= "000000";
      when 6253 => pixel <= "000000";
      when 6254 => pixel <= "000000";
      when 6255 => pixel <= "000000";
      when 6256 => pixel <= "000000";
      when 6257 => pixel <= "000000";
      when 6258 => pixel <= "000000";
      when 6259 => pixel <= "000000";
      when 6260 => pixel <= "000000";
      when 6261 => pixel <= "000000";
      when 6262 => pixel <= "000000";
      when 6263 => pixel <= "000000";
      when 6264 => pixel <= "000000";
      when 6265 => pixel <= "001101";
      when 6266 => pixel <= "001101";
      when 6267 => pixel <= "001101";
      when 6268 => pixel <= "001101";
      when 6269 => pixel <= "001101";
      when 6270 => pixel <= "001101";
      when 6271 => pixel <= "000000";
      when 6272 => pixel <= "000000";
      when 6273 => pixel <= "000000";
      when 6274 => pixel <= "001101";
      when 6275 => pixel <= "001101";
      when 6276 => pixel <= "001101";
      when 6277 => pixel <= "001101";
      when 6278 => pixel <= "001101";
      when 6279 => pixel <= "001101";
      when 6280 => pixel <= "000000";
      when 6281 => pixel <= "000000";
      when 6282 => pixel <= "000000";
      when 6283 => pixel <= "001101";
      when 6284 => pixel <= "001101";
      when 6285 => pixel <= "001101";
      when 6286 => pixel <= "001101";
      when 6287 => pixel <= "001101";
      when 6288 => pixel <= "001101";
      when 6289 => pixel <= "001101";
      when 6290 => pixel <= "000000";
      when 6291 => pixel <= "000000";
      when 6292 => pixel <= "000000";
      when 6293 => pixel <= "001101";
      when 6294 => pixel <= "001101";
      when 6295 => pixel <= "001101";
      when 6296 => pixel <= "001101";
      when 6297 => pixel <= "001101";
      when 6298 => pixel <= "000000";
      when 6299 => pixel <= "000000";
      when 6300 => pixel <= "000000";
      when 6301 => pixel <= "000000";
      when 6302 => pixel <= "001101";
      when 6303 => pixel <= "001101";
      when 6304 => pixel <= "001101";
      when 6305 => pixel <= "001101";
      when 6306 => pixel <= "001101";
      when 6307 => pixel <= "000000";
      when 6308 => pixel <= "000000";
      when 6309 => pixel <= "000000";
      when 6310 => pixel <= "000000";
      when 6311 => pixel <= "000000";
      when 6312 => pixel <= "000000";
      when 6313 => pixel <= "000000";
      when 6314 => pixel <= "000000";
      when 6315 => pixel <= "000000";
      when 6316 => pixel <= "000000";
      when 6317 => pixel <= "000000";
      when 6318 => pixel <= "000000";
      when 6319 => pixel <= "000000";
      when 6320 => pixel <= "000000";
      when 6321 => pixel <= "000000";
      when 6322 => pixel <= "000000";
      when 6323 => pixel <= "000000";
      when 6324 => pixel <= "001101";
      when 6325 => pixel <= "001101";
      when 6326 => pixel <= "000000";
      when 6327 => pixel <= "000000";
      when 6328 => pixel <= "000000";
      when 6329 => pixel <= "000000";
      when 6330 => pixel <= "000000";
      when 6331 => pixel <= "000000";
      when 6332 => pixel <= "001101";
      when 6333 => pixel <= "000000";
      when 6334 => pixel <= "000000";
      when 6335 => pixel <= "000000";
      when 6336 => pixel <= "000000";
      when 6337 => pixel <= "000000";
      when 6338 => pixel <= "000000";
      when 6339 => pixel <= "000000";
      when 6340 => pixel <= "001101";
      when 6341 => pixel <= "001101";
      when 6342 => pixel <= "000000";
      when 6343 => pixel <= "000000";
      when 6344 => pixel <= "000000";
      when 6345 => pixel <= "000000";
      when 6346 => pixel <= "000000";
      when 6347 => pixel <= "000000";
      when 6348 => pixel <= "000000";
      when 6349 => pixel <= "000000";
      when 6350 => pixel <= "000000";
      when 6351 => pixel <= "000000";
      when 6352 => pixel <= "000000";
      when 6353 => pixel <= "000000";
      when 6354 => pixel <= "000000";
      when 6355 => pixel <= "000000";
      when 6356 => pixel <= "000000";
      when 6357 => pixel <= "001101";
      when 6358 => pixel <= "001101";
      when 6359 => pixel <= "001101";
      when 6360 => pixel <= "001101";
      when 6361 => pixel <= "001101";
      when 6362 => pixel <= "001101";
      when 6363 => pixel <= "000000";
      when 6364 => pixel <= "000000";
      when 6365 => pixel <= "000000";
      when 6366 => pixel <= "001101";
      when 6367 => pixel <= "001101";
      when 6368 => pixel <= "001101";
      when 6369 => pixel <= "001101";
      when 6370 => pixel <= "001101";
      when 6371 => pixel <= "000000";
      when 6372 => pixel <= "000000";
      when 6373 => pixel <= "000000";
      when 6374 => pixel <= "000000";
      when 6375 => pixel <= "000000";
      when 6376 => pixel <= "000000";
      when 6377 => pixel <= "000000";
      when 6378 => pixel <= "000000";
      when 6379 => pixel <= "000000";
      when 6380 => pixel <= "000000";
      when 6381 => pixel <= "000000";
      when 6382 => pixel <= "000000";
      when 6383 => pixel <= "000000";
      when 6384 => pixel <= "000000";
      when 6385 => pixel <= "000000";
      when 6386 => pixel <= "000000";
      when 6387 => pixel <= "000000";
      when 6388 => pixel <= "000000";
      when 6389 => pixel <= "000000";
      when 6390 => pixel <= "000000";
      when 6391 => pixel <= "000000";
      when 6392 => pixel <= "000000";
      when 6393 => pixel <= "000000";
      when 6394 => pixel <= "000000";
      when 6395 => pixel <= "000000";
      when 6396 => pixel <= "000000";
      when 6397 => pixel <= "000000";
      when 6398 => pixel <= "000000";
      when 6399 => pixel <= "000000";
      when 6400 => pixel <= "000000";
      when 6401 => pixel <= "000000";
      when 6402 => pixel <= "000000";
      when 6403 => pixel <= "000000";
      when 6404 => pixel <= "000000";
      when 6405 => pixel <= "000000";
      when 6406 => pixel <= "000000";
      when 6407 => pixel <= "000000";
      when 6408 => pixel <= "000000";
      when 6409 => pixel <= "000000";
      when 6410 => pixel <= "000000";
      when 6411 => pixel <= "000000";
      when 6412 => pixel <= "000000";
      when 6413 => pixel <= "000000";
      when 6414 => pixel <= "000000";
      when 6415 => pixel <= "000000";
      when 6416 => pixel <= "000000";
      when 6417 => pixel <= "000000";
      when 6418 => pixel <= "000000";
      when 6419 => pixel <= "000000";
      when 6420 => pixel <= "000000";
      when 6421 => pixel <= "000000";
      when 6422 => pixel <= "000000";
      when 6423 => pixel <= "000000";
      when 6424 => pixel <= "000000";
      when 6425 => pixel <= "000000";
      when 6426 => pixel <= "001101";
      when 6427 => pixel <= "001101";
      when 6428 => pixel <= "000000";
      when 6429 => pixel <= "000000";
      when 6430 => pixel <= "001101";
      when 6431 => pixel <= "001101";
      when 6432 => pixel <= "000000";
      when 6433 => pixel <= "000000";
      when 6434 => pixel <= "000000";
      when 6435 => pixel <= "001101";
      when 6436 => pixel <= "001101";
      when 6437 => pixel <= "000000";
      when 6438 => pixel <= "000000";
      when 6439 => pixel <= "001101";
      when 6440 => pixel <= "001101";
      when 6441 => pixel <= "000000";
      when 6442 => pixel <= "000000";
      when 6443 => pixel <= "000000";
      when 6444 => pixel <= "001101";
      when 6445 => pixel <= "001101";
      when 6446 => pixel <= "000000";
      when 6447 => pixel <= "000000";
      when 6448 => pixel <= "001101";
      when 6449 => pixel <= "001101";
      when 6450 => pixel <= "000000";
      when 6451 => pixel <= "000000";
      when 6452 => pixel <= "001101";
      when 6453 => pixel <= "001101";
      when 6454 => pixel <= "000000";
      when 6455 => pixel <= "000000";
      when 6456 => pixel <= "000000";
      when 6457 => pixel <= "001101";
      when 6458 => pixel <= "001101";
      when 6459 => pixel <= "000000";
      when 6460 => pixel <= "000000";
      when 6461 => pixel <= "001101";
      when 6462 => pixel <= "001101";
      when 6463 => pixel <= "000000";
      when 6464 => pixel <= "000000";
      when 6465 => pixel <= "000000";
      when 6466 => pixel <= "001101";
      when 6467 => pixel <= "001101";
      when 6468 => pixel <= "000000";
      when 6469 => pixel <= "000000";
      when 6470 => pixel <= "000000";
      when 6471 => pixel <= "000000";
      when 6472 => pixel <= "000000";
      when 6473 => pixel <= "000000";
      when 6474 => pixel <= "000000";
      when 6475 => pixel <= "000000";
      when 6476 => pixel <= "000000";
      when 6477 => pixel <= "000000";
      when 6478 => pixel <= "000000";
      when 6479 => pixel <= "000000";
      when 6480 => pixel <= "000000";
      when 6481 => pixel <= "000000";
      when 6482 => pixel <= "000000";
      when 6483 => pixel <= "001101";
      when 6484 => pixel <= "001101";
      when 6485 => pixel <= "000000";
      when 6486 => pixel <= "000000";
      when 6487 => pixel <= "000000";
      when 6488 => pixel <= "000000";
      when 6489 => pixel <= "000000";
      when 6490 => pixel <= "000000";
      when 6491 => pixel <= "001101";
      when 6492 => pixel <= "001101";
      when 6493 => pixel <= "001101";
      when 6494 => pixel <= "000000";
      when 6495 => pixel <= "000000";
      when 6496 => pixel <= "000000";
      when 6497 => pixel <= "000000";
      when 6498 => pixel <= "000000";
      when 6499 => pixel <= "000000";
      when 6500 => pixel <= "000000";
      when 6501 => pixel <= "001101";
      when 6502 => pixel <= "001101";
      when 6503 => pixel <= "000000";
      when 6504 => pixel <= "000000";
      when 6505 => pixel <= "000000";
      when 6506 => pixel <= "000000";
      when 6507 => pixel <= "000000";
      when 6508 => pixel <= "000000";
      when 6509 => pixel <= "000000";
      when 6510 => pixel <= "000000";
      when 6511 => pixel <= "000000";
      when 6512 => pixel <= "000000";
      when 6513 => pixel <= "000000";
      when 6514 => pixel <= "000000";
      when 6515 => pixel <= "000000";
      when 6516 => pixel <= "000000";
      when 6517 => pixel <= "001101";
      when 6518 => pixel <= "001101";
      when 6519 => pixel <= "001101";
      when 6520 => pixel <= "001101";
      when 6521 => pixel <= "001101";
      when 6522 => pixel <= "001101";
      when 6523 => pixel <= "000000";
      when 6524 => pixel <= "000000";
      when 6525 => pixel <= "001101";
      when 6526 => pixel <= "001101";
      when 6527 => pixel <= "000000";
      when 6528 => pixel <= "000000";
      when 6529 => pixel <= "000000";
      when 6530 => pixel <= "001101";
      when 6531 => pixel <= "001101";
      when 6532 => pixel <= "000000";
      when 6533 => pixel <= "000000";
      when 6534 => pixel <= "000000";
      when 6535 => pixel <= "000000";
      when 6536 => pixel <= "000000";
      when 6537 => pixel <= "000000";
      when 6538 => pixel <= "000000";
      when 6539 => pixel <= "000000";
      when 6540 => pixel <= "000000";
      when 6541 => pixel <= "000000";
      when 6542 => pixel <= "000000";
      when 6543 => pixel <= "000000";
      when 6544 => pixel <= "000000";
      when 6545 => pixel <= "000000";
      when 6546 => pixel <= "000000";
      when 6547 => pixel <= "000000";
      when 6548 => pixel <= "000000";
      when 6549 => pixel <= "000000";
      when 6550 => pixel <= "000000";
      when 6551 => pixel <= "000000";
      when 6552 => pixel <= "000000";
      when 6553 => pixel <= "000000";
      when 6554 => pixel <= "000000";
      when 6555 => pixel <= "000000";
      when 6556 => pixel <= "000000";
      when 6557 => pixel <= "000000";
      when 6558 => pixel <= "000000";
      when 6559 => pixel <= "000000";
      when 6560 => pixel <= "000000";
      when 6561 => pixel <= "000000";
      when 6562 => pixel <= "000000";
      when 6563 => pixel <= "000000";
      when 6564 => pixel <= "000000";
      when 6565 => pixel <= "000000";
      when 6566 => pixel <= "000000";
      when 6567 => pixel <= "000000";
      when 6568 => pixel <= "000000";
      when 6569 => pixel <= "000000";
      when 6570 => pixel <= "000000";
      when 6571 => pixel <= "000000";
      when 6572 => pixel <= "000000";
      when 6573 => pixel <= "000000";
      when 6574 => pixel <= "000000";
      when 6575 => pixel <= "000000";
      when 6576 => pixel <= "000000";
      when 6577 => pixel <= "000000";
      when 6578 => pixel <= "000000";
      when 6579 => pixel <= "000000";
      when 6580 => pixel <= "000000";
      when 6581 => pixel <= "000000";
      when 6582 => pixel <= "000000";
      when 6583 => pixel <= "000000";
      when 6584 => pixel <= "000000";
      when 6585 => pixel <= "000000";
      when 6586 => pixel <= "001101";
      when 6587 => pixel <= "001101";
      when 6588 => pixel <= "000000";
      when 6589 => pixel <= "000000";
      when 6590 => pixel <= "001101";
      when 6591 => pixel <= "001101";
      when 6592 => pixel <= "000000";
      when 6593 => pixel <= "000000";
      when 6594 => pixel <= "000000";
      when 6595 => pixel <= "001101";
      when 6596 => pixel <= "001101";
      when 6597 => pixel <= "000000";
      when 6598 => pixel <= "000000";
      when 6599 => pixel <= "001101";
      when 6600 => pixel <= "001101";
      when 6601 => pixel <= "000000";
      when 6602 => pixel <= "000000";
      when 6603 => pixel <= "000000";
      when 6604 => pixel <= "001101";
      when 6605 => pixel <= "001101";
      when 6606 => pixel <= "000000";
      when 6607 => pixel <= "000000";
      when 6608 => pixel <= "000000";
      when 6609 => pixel <= "001101";
      when 6610 => pixel <= "000000";
      when 6611 => pixel <= "000000";
      when 6612 => pixel <= "001101";
      when 6613 => pixel <= "001101";
      when 6614 => pixel <= "000000";
      when 6615 => pixel <= "000000";
      when 6616 => pixel <= "000000";
      when 6617 => pixel <= "001101";
      when 6618 => pixel <= "001101";
      when 6619 => pixel <= "000000";
      when 6620 => pixel <= "000000";
      when 6621 => pixel <= "001101";
      when 6622 => pixel <= "001101";
      when 6623 => pixel <= "000000";
      when 6624 => pixel <= "000000";
      when 6625 => pixel <= "000000";
      when 6626 => pixel <= "001101";
      when 6627 => pixel <= "001101";
      when 6628 => pixel <= "000000";
      when 6629 => pixel <= "000000";
      when 6630 => pixel <= "000000";
      when 6631 => pixel <= "000000";
      when 6632 => pixel <= "000000";
      when 6633 => pixel <= "000000";
      when 6634 => pixel <= "000000";
      when 6635 => pixel <= "000000";
      when 6636 => pixel <= "000000";
      when 6637 => pixel <= "000000";
      when 6638 => pixel <= "000000";
      when 6639 => pixel <= "000000";
      when 6640 => pixel <= "000000";
      when 6641 => pixel <= "000000";
      when 6642 => pixel <= "001101";
      when 6643 => pixel <= "001101";
      when 6644 => pixel <= "000000";
      when 6645 => pixel <= "000000";
      when 6646 => pixel <= "000000";
      when 6647 => pixel <= "000000";
      when 6648 => pixel <= "000000";
      when 6649 => pixel <= "000000";
      when 6650 => pixel <= "001101";
      when 6651 => pixel <= "001101";
      when 6652 => pixel <= "000000";
      when 6653 => pixel <= "001101";
      when 6654 => pixel <= "001101";
      when 6655 => pixel <= "000000";
      when 6656 => pixel <= "000000";
      when 6657 => pixel <= "000000";
      when 6658 => pixel <= "000000";
      when 6659 => pixel <= "000000";
      when 6660 => pixel <= "000000";
      when 6661 => pixel <= "000000";
      when 6662 => pixel <= "001101";
      when 6663 => pixel <= "001101";
      when 6664 => pixel <= "000000";
      when 6665 => pixel <= "000000";
      when 6666 => pixel <= "000000";
      when 6667 => pixel <= "000000";
      when 6668 => pixel <= "000000";
      when 6669 => pixel <= "000000";
      when 6670 => pixel <= "000000";
      when 6671 => pixel <= "000000";
      when 6672 => pixel <= "000000";
      when 6673 => pixel <= "000000";
      when 6674 => pixel <= "000000";
      when 6675 => pixel <= "000000";
      when 6676 => pixel <= "000000";
      when 6677 => pixel <= "001101";
      when 6678 => pixel <= "000000";
      when 6679 => pixel <= "001101";
      when 6680 => pixel <= "001101";
      when 6681 => pixel <= "000000";
      when 6682 => pixel <= "001101";
      when 6683 => pixel <= "000000";
      when 6684 => pixel <= "000000";
      when 6685 => pixel <= "001101";
      when 6686 => pixel <= "001101";
      when 6687 => pixel <= "000000";
      when 6688 => pixel <= "000000";
      when 6689 => pixel <= "000000";
      when 6690 => pixel <= "001101";
      when 6691 => pixel <= "001101";
      when 6692 => pixel <= "000000";
      when 6693 => pixel <= "000000";
      when 6694 => pixel <= "000000";
      when 6695 => pixel <= "000000";
      when 6696 => pixel <= "000000";
      when 6697 => pixel <= "000000";
      when 6698 => pixel <= "000000";
      when 6699 => pixel <= "000000";
      when 6700 => pixel <= "000000";
      when 6701 => pixel <= "000000";
      when 6702 => pixel <= "000000";
      when 6703 => pixel <= "000000";
      when 6704 => pixel <= "000000";
      when 6705 => pixel <= "000000";
      when 6706 => pixel <= "000000";
      when 6707 => pixel <= "000000";
      when 6708 => pixel <= "000000";
      when 6709 => pixel <= "000000";
      when 6710 => pixel <= "000000";
      when 6711 => pixel <= "000000";
      when 6712 => pixel <= "000000";
      when 6713 => pixel <= "000000";
      when 6714 => pixel <= "000000";
      when 6715 => pixel <= "000000";
      when 6716 => pixel <= "000000";
      when 6717 => pixel <= "000000";
      when 6718 => pixel <= "000000";
      when 6719 => pixel <= "000000";
      when 6720 => pixel <= "000000";
      when 6721 => pixel <= "000000";
      when 6722 => pixel <= "000000";
      when 6723 => pixel <= "000000";
      when 6724 => pixel <= "000000";
      when 6725 => pixel <= "000000";
      when 6726 => pixel <= "000000";
      when 6727 => pixel <= "000000";
      when 6728 => pixel <= "000000";
      when 6729 => pixel <= "000000";
      when 6730 => pixel <= "000000";
      when 6731 => pixel <= "000000";
      when 6732 => pixel <= "000000";
      when 6733 => pixel <= "000000";
      when 6734 => pixel <= "000000";
      when 6735 => pixel <= "000000";
      when 6736 => pixel <= "000000";
      when 6737 => pixel <= "000000";
      when 6738 => pixel <= "000000";
      when 6739 => pixel <= "000000";
      when 6740 => pixel <= "000000";
      when 6741 => pixel <= "000000";
      when 6742 => pixel <= "000000";
      when 6743 => pixel <= "000000";
      when 6744 => pixel <= "000000";
      when 6745 => pixel <= "000000";
      when 6746 => pixel <= "001101";
      when 6747 => pixel <= "001101";
      when 6748 => pixel <= "000000";
      when 6749 => pixel <= "000000";
      when 6750 => pixel <= "001101";
      when 6751 => pixel <= "001101";
      when 6752 => pixel <= "000000";
      when 6753 => pixel <= "000000";
      when 6754 => pixel <= "000000";
      when 6755 => pixel <= "001101";
      when 6756 => pixel <= "001101";
      when 6757 => pixel <= "000000";
      when 6758 => pixel <= "000000";
      when 6759 => pixel <= "001101";
      when 6760 => pixel <= "001101";
      when 6761 => pixel <= "000000";
      when 6762 => pixel <= "000000";
      when 6763 => pixel <= "000000";
      when 6764 => pixel <= "001101";
      when 6765 => pixel <= "001101";
      when 6766 => pixel <= "000000";
      when 6767 => pixel <= "001101";
      when 6768 => pixel <= "000000";
      when 6769 => pixel <= "000000";
      when 6770 => pixel <= "000000";
      when 6771 => pixel <= "000000";
      when 6772 => pixel <= "000000";
      when 6773 => pixel <= "001101";
      when 6774 => pixel <= "001101";
      when 6775 => pixel <= "000000";
      when 6776 => pixel <= "000000";
      when 6777 => pixel <= "000000";
      when 6778 => pixel <= "000000";
      when 6779 => pixel <= "000000";
      when 6780 => pixel <= "000000";
      when 6781 => pixel <= "000000";
      when 6782 => pixel <= "001101";
      when 6783 => pixel <= "001101";
      when 6784 => pixel <= "000000";
      when 6785 => pixel <= "000000";
      when 6786 => pixel <= "000000";
      when 6787 => pixel <= "000000";
      when 6788 => pixel <= "000000";
      when 6789 => pixel <= "000000";
      when 6790 => pixel <= "000000";
      when 6791 => pixel <= "000000";
      when 6792 => pixel <= "000000";
      when 6793 => pixel <= "000000";
      when 6794 => pixel <= "000000";
      when 6795 => pixel <= "000000";
      when 6796 => pixel <= "000000";
      when 6797 => pixel <= "000000";
      when 6798 => pixel <= "000000";
      when 6799 => pixel <= "000000";
      when 6800 => pixel <= "000000";
      when 6801 => pixel <= "000000";
      when 6802 => pixel <= "001101";
      when 6803 => pixel <= "001101";
      when 6804 => pixel <= "000000";
      when 6805 => pixel <= "000000";
      when 6806 => pixel <= "000000";
      when 6807 => pixel <= "000000";
      when 6808 => pixel <= "000000";
      when 6809 => pixel <= "001101";
      when 6810 => pixel <= "001101";
      when 6811 => pixel <= "000000";
      when 6812 => pixel <= "000000";
      when 6813 => pixel <= "000000";
      when 6814 => pixel <= "001101";
      when 6815 => pixel <= "001101";
      when 6816 => pixel <= "000000";
      when 6817 => pixel <= "000000";
      when 6818 => pixel <= "000000";
      when 6819 => pixel <= "000000";
      when 6820 => pixel <= "000000";
      when 6821 => pixel <= "000000";
      when 6822 => pixel <= "001101";
      when 6823 => pixel <= "001101";
      when 6824 => pixel <= "000000";
      when 6825 => pixel <= "000000";
      when 6826 => pixel <= "000000";
      when 6827 => pixel <= "000000";
      when 6828 => pixel <= "000000";
      when 6829 => pixel <= "000000";
      when 6830 => pixel <= "000000";
      when 6831 => pixel <= "000000";
      when 6832 => pixel <= "000000";
      when 6833 => pixel <= "000000";
      when 6834 => pixel <= "000000";
      when 6835 => pixel <= "000000";
      when 6836 => pixel <= "000000";
      when 6837 => pixel <= "000000";
      when 6838 => pixel <= "000000";
      when 6839 => pixel <= "001101";
      when 6840 => pixel <= "001101";
      when 6841 => pixel <= "000000";
      when 6842 => pixel <= "000000";
      when 6843 => pixel <= "000000";
      when 6844 => pixel <= "000000";
      when 6845 => pixel <= "001101";
      when 6846 => pixel <= "001101";
      when 6847 => pixel <= "000000";
      when 6848 => pixel <= "000000";
      when 6849 => pixel <= "000000";
      when 6850 => pixel <= "001101";
      when 6851 => pixel <= "001101";
      when 6852 => pixel <= "000000";
      when 6853 => pixel <= "000000";
      when 6854 => pixel <= "000000";
      when 6855 => pixel <= "000000";
      when 6856 => pixel <= "000000";
      when 6857 => pixel <= "000000";
      when 6858 => pixel <= "000000";
      when 6859 => pixel <= "000000";
      when 6860 => pixel <= "000000";
      when 6861 => pixel <= "000000";
      when 6862 => pixel <= "000000";
      when 6863 => pixel <= "000000";
      when 6864 => pixel <= "000000";
      when 6865 => pixel <= "000000";
      when 6866 => pixel <= "000000";
      when 6867 => pixel <= "000000";
      when 6868 => pixel <= "000000";
      when 6869 => pixel <= "000000";
      when 6870 => pixel <= "000000";
      when 6871 => pixel <= "000000";
      when 6872 => pixel <= "000000";
      when 6873 => pixel <= "000000";
      when 6874 => pixel <= "000000";
      when 6875 => pixel <= "000000";
      when 6876 => pixel <= "000000";
      when 6877 => pixel <= "000000";
      when 6878 => pixel <= "000000";
      when 6879 => pixel <= "000000";
      when 6880 => pixel <= "000000";
      when 6881 => pixel <= "000000";
      when 6882 => pixel <= "000000";
      when 6883 => pixel <= "000000";
      when 6884 => pixel <= "000000";
      when 6885 => pixel <= "000000";
      when 6886 => pixel <= "000000";
      when 6887 => pixel <= "000000";
      when 6888 => pixel <= "000000";
      when 6889 => pixel <= "000000";
      when 6890 => pixel <= "000000";
      when 6891 => pixel <= "000000";
      when 6892 => pixel <= "000000";
      when 6893 => pixel <= "000000";
      when 6894 => pixel <= "000000";
      when 6895 => pixel <= "000000";
      when 6896 => pixel <= "000000";
      when 6897 => pixel <= "000000";
      when 6898 => pixel <= "000000";
      when 6899 => pixel <= "000000";
      when 6900 => pixel <= "000000";
      when 6901 => pixel <= "000000";
      when 6902 => pixel <= "000000";
      when 6903 => pixel <= "000000";
      when 6904 => pixel <= "000000";
      when 6905 => pixel <= "000000";
      when 6906 => pixel <= "001101";
      when 6907 => pixel <= "001101";
      when 6908 => pixel <= "001101";
      when 6909 => pixel <= "001101";
      when 6910 => pixel <= "001101";
      when 6911 => pixel <= "000000";
      when 6912 => pixel <= "000000";
      when 6913 => pixel <= "000000";
      when 6914 => pixel <= "000000";
      when 6915 => pixel <= "001101";
      when 6916 => pixel <= "001101";
      when 6917 => pixel <= "001101";
      when 6918 => pixel <= "001101";
      when 6919 => pixel <= "001101";
      when 6920 => pixel <= "000000";
      when 6921 => pixel <= "000000";
      when 6922 => pixel <= "000000";
      when 6923 => pixel <= "000000";
      when 6924 => pixel <= "001101";
      when 6925 => pixel <= "001101";
      when 6926 => pixel <= "001101";
      when 6927 => pixel <= "001101";
      when 6928 => pixel <= "000000";
      when 6929 => pixel <= "000000";
      when 6930 => pixel <= "000000";
      when 6931 => pixel <= "000000";
      when 6932 => pixel <= "000000";
      when 6933 => pixel <= "000000";
      when 6934 => pixel <= "001101";
      when 6935 => pixel <= "001101";
      when 6936 => pixel <= "001101";
      when 6937 => pixel <= "000000";
      when 6938 => pixel <= "000000";
      when 6939 => pixel <= "000000";
      when 6940 => pixel <= "000000";
      when 6941 => pixel <= "000000";
      when 6942 => pixel <= "000000";
      when 6943 => pixel <= "001101";
      when 6944 => pixel <= "001101";
      when 6945 => pixel <= "001101";
      when 6946 => pixel <= "000000";
      when 6947 => pixel <= "000000";
      when 6948 => pixel <= "000000";
      when 6949 => pixel <= "000000";
      when 6950 => pixel <= "000000";
      when 6951 => pixel <= "000000";
      when 6952 => pixel <= "000000";
      when 6953 => pixel <= "000000";
      when 6954 => pixel <= "000000";
      when 6955 => pixel <= "000000";
      when 6956 => pixel <= "000000";
      when 6957 => pixel <= "000000";
      when 6958 => pixel <= "000000";
      when 6959 => pixel <= "000000";
      when 6960 => pixel <= "000000";
      when 6961 => pixel <= "000000";
      when 6962 => pixel <= "001101";
      when 6963 => pixel <= "001101";
      when 6964 => pixel <= "000000";
      when 6965 => pixel <= "000000";
      when 6966 => pixel <= "000000";
      when 6967 => pixel <= "000000";
      when 6968 => pixel <= "000000";
      when 6969 => pixel <= "001101";
      when 6970 => pixel <= "001101";
      when 6971 => pixel <= "000000";
      when 6972 => pixel <= "000000";
      when 6973 => pixel <= "000000";
      when 6974 => pixel <= "001101";
      when 6975 => pixel <= "001101";
      when 6976 => pixel <= "000000";
      when 6977 => pixel <= "000000";
      when 6978 => pixel <= "000000";
      when 6979 => pixel <= "000000";
      when 6980 => pixel <= "000000";
      when 6981 => pixel <= "000000";
      when 6982 => pixel <= "001101";
      when 6983 => pixel <= "001101";
      when 6984 => pixel <= "000000";
      when 6985 => pixel <= "000000";
      when 6986 => pixel <= "000000";
      when 6987 => pixel <= "000000";
      when 6988 => pixel <= "000000";
      when 6989 => pixel <= "000000";
      when 6990 => pixel <= "000000";
      when 6991 => pixel <= "000000";
      when 6992 => pixel <= "000000";
      when 6993 => pixel <= "000000";
      when 6994 => pixel <= "000000";
      when 6995 => pixel <= "000000";
      when 6996 => pixel <= "000000";
      when 6997 => pixel <= "000000";
      when 6998 => pixel <= "000000";
      when 6999 => pixel <= "001101";
      when 7000 => pixel <= "001101";
      when 7001 => pixel <= "000000";
      when 7002 => pixel <= "000000";
      when 7003 => pixel <= "000000";
      when 7004 => pixel <= "000000";
      when 7005 => pixel <= "001101";
      when 7006 => pixel <= "001101";
      when 7007 => pixel <= "000000";
      when 7008 => pixel <= "000000";
      when 7009 => pixel <= "000000";
      when 7010 => pixel <= "001101";
      when 7011 => pixel <= "001101";
      when 7012 => pixel <= "000000";
      when 7013 => pixel <= "000000";
      when 7014 => pixel <= "000000";
      when 7015 => pixel <= "000000";
      when 7016 => pixel <= "000000";
      when 7017 => pixel <= "000000";
      when 7018 => pixel <= "000000";
      when 7019 => pixel <= "000000";
      when 7020 => pixel <= "000000";
      when 7021 => pixel <= "000000";
      when 7022 => pixel <= "000000";
      when 7023 => pixel <= "000000";
      when 7024 => pixel <= "000000";
      when 7025 => pixel <= "000000";
      when 7026 => pixel <= "000000";
      when 7027 => pixel <= "000000";
      when 7028 => pixel <= "000000";
      when 7029 => pixel <= "000000";
      when 7030 => pixel <= "000000";
      when 7031 => pixel <= "000000";
      when 7032 => pixel <= "000000";
      when 7033 => pixel <= "000000";
      when 7034 => pixel <= "000000";
      when 7035 => pixel <= "000000";
      when 7036 => pixel <= "000000";
      when 7037 => pixel <= "000000";
      when 7038 => pixel <= "000000";
      when 7039 => pixel <= "000000";
      when 7040 => pixel <= "000000";
      when 7041 => pixel <= "000000";
      when 7042 => pixel <= "000000";
      when 7043 => pixel <= "000000";
      when 7044 => pixel <= "000000";
      when 7045 => pixel <= "000000";
      when 7046 => pixel <= "000000";
      when 7047 => pixel <= "000000";
      when 7048 => pixel <= "000000";
      when 7049 => pixel <= "000000";
      when 7050 => pixel <= "000000";
      when 7051 => pixel <= "000000";
      when 7052 => pixel <= "000000";
      when 7053 => pixel <= "000000";
      when 7054 => pixel <= "000000";
      when 7055 => pixel <= "000000";
      when 7056 => pixel <= "000000";
      when 7057 => pixel <= "000000";
      when 7058 => pixel <= "000000";
      when 7059 => pixel <= "000000";
      when 7060 => pixel <= "000000";
      when 7061 => pixel <= "000000";
      when 7062 => pixel <= "000000";
      when 7063 => pixel <= "000000";
      when 7064 => pixel <= "000000";
      when 7065 => pixel <= "000000";
      when 7066 => pixel <= "001101";
      when 7067 => pixel <= "001101";
      when 7068 => pixel <= "000000";
      when 7069 => pixel <= "000000";
      when 7070 => pixel <= "000000";
      when 7071 => pixel <= "000000";
      when 7072 => pixel <= "000000";
      when 7073 => pixel <= "000000";
      when 7074 => pixel <= "000000";
      when 7075 => pixel <= "001101";
      when 7076 => pixel <= "001101";
      when 7077 => pixel <= "000000";
      when 7078 => pixel <= "001101";
      when 7079 => pixel <= "001101";
      when 7080 => pixel <= "000000";
      when 7081 => pixel <= "000000";
      when 7082 => pixel <= "000000";
      when 7083 => pixel <= "000000";
      when 7084 => pixel <= "001101";
      when 7085 => pixel <= "001101";
      when 7086 => pixel <= "000000";
      when 7087 => pixel <= "001101";
      when 7088 => pixel <= "000000";
      when 7089 => pixel <= "000000";
      when 7090 => pixel <= "000000";
      when 7091 => pixel <= "000000";
      when 7092 => pixel <= "000000";
      when 7093 => pixel <= "000000";
      when 7094 => pixel <= "000000";
      when 7095 => pixel <= "000000";
      when 7096 => pixel <= "001101";
      when 7097 => pixel <= "001101";
      when 7098 => pixel <= "000000";
      when 7099 => pixel <= "000000";
      when 7100 => pixel <= "000000";
      when 7101 => pixel <= "000000";
      when 7102 => pixel <= "000000";
      when 7103 => pixel <= "000000";
      when 7104 => pixel <= "000000";
      when 7105 => pixel <= "001101";
      when 7106 => pixel <= "001101";
      when 7107 => pixel <= "000000";
      when 7108 => pixel <= "000000";
      when 7109 => pixel <= "000000";
      when 7110 => pixel <= "000000";
      when 7111 => pixel <= "000000";
      when 7112 => pixel <= "000000";
      when 7113 => pixel <= "000000";
      when 7114 => pixel <= "000000";
      when 7115 => pixel <= "000000";
      when 7116 => pixel <= "000000";
      when 7117 => pixel <= "000000";
      when 7118 => pixel <= "000000";
      when 7119 => pixel <= "000000";
      when 7120 => pixel <= "000000";
      when 7121 => pixel <= "000000";
      when 7122 => pixel <= "001101";
      when 7123 => pixel <= "001101";
      when 7124 => pixel <= "000000";
      when 7125 => pixel <= "000000";
      when 7126 => pixel <= "000000";
      when 7127 => pixel <= "000000";
      when 7128 => pixel <= "000000";
      when 7129 => pixel <= "001101";
      when 7130 => pixel <= "001101";
      when 7131 => pixel <= "001101";
      when 7132 => pixel <= "001101";
      when 7133 => pixel <= "001101";
      when 7134 => pixel <= "001101";
      when 7135 => pixel <= "001101";
      when 7136 => pixel <= "000000";
      when 7137 => pixel <= "000000";
      when 7138 => pixel <= "000000";
      when 7139 => pixel <= "000000";
      when 7140 => pixel <= "000000";
      when 7141 => pixel <= "000000";
      when 7142 => pixel <= "001101";
      when 7143 => pixel <= "001101";
      when 7144 => pixel <= "000000";
      when 7145 => pixel <= "000000";
      when 7146 => pixel <= "000000";
      when 7147 => pixel <= "000000";
      when 7148 => pixel <= "000000";
      when 7149 => pixel <= "000000";
      when 7150 => pixel <= "000000";
      when 7151 => pixel <= "000000";
      when 7152 => pixel <= "000000";
      when 7153 => pixel <= "000000";
      when 7154 => pixel <= "000000";
      when 7155 => pixel <= "000000";
      when 7156 => pixel <= "000000";
      when 7157 => pixel <= "000000";
      when 7158 => pixel <= "000000";
      when 7159 => pixel <= "001101";
      when 7160 => pixel <= "001101";
      when 7161 => pixel <= "000000";
      when 7162 => pixel <= "000000";
      when 7163 => pixel <= "000000";
      when 7164 => pixel <= "000000";
      when 7165 => pixel <= "001101";
      when 7166 => pixel <= "001101";
      when 7167 => pixel <= "000000";
      when 7168 => pixel <= "000000";
      when 7169 => pixel <= "000000";
      when 7170 => pixel <= "001101";
      when 7171 => pixel <= "001101";
      when 7172 => pixel <= "000000";
      when 7173 => pixel <= "000000";
      when 7174 => pixel <= "000000";
      when 7175 => pixel <= "000000";
      when 7176 => pixel <= "000000";
      when 7177 => pixel <= "000000";
      when 7178 => pixel <= "000000";
      when 7179 => pixel <= "000000";
      when 7180 => pixel <= "000000";
      when 7181 => pixel <= "000000";
      when 7182 => pixel <= "000000";
      when 7183 => pixel <= "000000";
      when 7184 => pixel <= "000000";
      when 7185 => pixel <= "000000";
      when 7186 => pixel <= "000000";
      when 7187 => pixel <= "000000";
      when 7188 => pixel <= "000000";
      when 7189 => pixel <= "000000";
      when 7190 => pixel <= "000000";
      when 7191 => pixel <= "000000";
      when 7192 => pixel <= "000000";
      when 7193 => pixel <= "000000";
      when 7194 => pixel <= "000000";
      when 7195 => pixel <= "000000";
      when 7196 => pixel <= "000000";
      when 7197 => pixel <= "000000";
      when 7198 => pixel <= "000000";
      when 7199 => pixel <= "000000";
      when 7200 => pixel <= "000000";
      when 7201 => pixel <= "000000";
      when 7202 => pixel <= "000000";
      when 7203 => pixel <= "000000";
      when 7204 => pixel <= "000000";
      when 7205 => pixel <= "000000";
      when 7206 => pixel <= "000000";
      when 7207 => pixel <= "000000";
      when 7208 => pixel <= "000000";
      when 7209 => pixel <= "000000";
      when 7210 => pixel <= "000000";
      when 7211 => pixel <= "000000";
      when 7212 => pixel <= "000000";
      when 7213 => pixel <= "000000";
      when 7214 => pixel <= "000000";
      when 7215 => pixel <= "000000";
      when 7216 => pixel <= "000000";
      when 7217 => pixel <= "000000";
      when 7218 => pixel <= "000000";
      when 7219 => pixel <= "000000";
      when 7220 => pixel <= "000000";
      when 7221 => pixel <= "000000";
      when 7222 => pixel <= "000000";
      when 7223 => pixel <= "000000";
      when 7224 => pixel <= "000000";
      when 7225 => pixel <= "000000";
      when 7226 => pixel <= "001101";
      when 7227 => pixel <= "001101";
      when 7228 => pixel <= "000000";
      when 7229 => pixel <= "000000";
      when 7230 => pixel <= "000000";
      when 7231 => pixel <= "000000";
      when 7232 => pixel <= "000000";
      when 7233 => pixel <= "000000";
      when 7234 => pixel <= "000000";
      when 7235 => pixel <= "001101";
      when 7236 => pixel <= "001101";
      when 7237 => pixel <= "000000";
      when 7238 => pixel <= "000000";
      when 7239 => pixel <= "001101";
      when 7240 => pixel <= "001101";
      when 7241 => pixel <= "000000";
      when 7242 => pixel <= "000000";
      when 7243 => pixel <= "000000";
      when 7244 => pixel <= "001101";
      when 7245 => pixel <= "001101";
      when 7246 => pixel <= "000000";
      when 7247 => pixel <= "000000";
      when 7248 => pixel <= "000000";
      when 7249 => pixel <= "000000";
      when 7250 => pixel <= "000000";
      when 7251 => pixel <= "000000";
      when 7252 => pixel <= "000000";
      when 7253 => pixel <= "000000";
      when 7254 => pixel <= "000000";
      when 7255 => pixel <= "000000";
      when 7256 => pixel <= "000000";
      when 7257 => pixel <= "001101";
      when 7258 => pixel <= "001101";
      when 7259 => pixel <= "000000";
      when 7260 => pixel <= "000000";
      when 7261 => pixel <= "000000";
      when 7262 => pixel <= "000000";
      when 7263 => pixel <= "000000";
      when 7264 => pixel <= "000000";
      when 7265 => pixel <= "000000";
      when 7266 => pixel <= "001101";
      when 7267 => pixel <= "001101";
      when 7268 => pixel <= "000000";
      when 7269 => pixel <= "000000";
      when 7270 => pixel <= "000000";
      when 7271 => pixel <= "000000";
      when 7272 => pixel <= "000000";
      when 7273 => pixel <= "000000";
      when 7274 => pixel <= "000000";
      when 7275 => pixel <= "000000";
      when 7276 => pixel <= "000000";
      when 7277 => pixel <= "000000";
      when 7278 => pixel <= "000000";
      when 7279 => pixel <= "000000";
      when 7280 => pixel <= "000000";
      when 7281 => pixel <= "000000";
      when 7282 => pixel <= "001101";
      when 7283 => pixel <= "001101";
      when 7284 => pixel <= "000000";
      when 7285 => pixel <= "000000";
      when 7286 => pixel <= "000000";
      when 7287 => pixel <= "000000";
      when 7288 => pixel <= "000000";
      when 7289 => pixel <= "001101";
      when 7290 => pixel <= "001101";
      when 7291 => pixel <= "000000";
      when 7292 => pixel <= "000000";
      when 7293 => pixel <= "000000";
      when 7294 => pixel <= "001101";
      when 7295 => pixel <= "001101";
      when 7296 => pixel <= "000000";
      when 7297 => pixel <= "000000";
      when 7298 => pixel <= "000000";
      when 7299 => pixel <= "000000";
      when 7300 => pixel <= "000000";
      when 7301 => pixel <= "000000";
      when 7302 => pixel <= "001101";
      when 7303 => pixel <= "001101";
      when 7304 => pixel <= "000000";
      when 7305 => pixel <= "000000";
      when 7306 => pixel <= "000000";
      when 7307 => pixel <= "000000";
      when 7308 => pixel <= "000000";
      when 7309 => pixel <= "000000";
      when 7310 => pixel <= "000000";
      when 7311 => pixel <= "000000";
      when 7312 => pixel <= "000000";
      when 7313 => pixel <= "000000";
      when 7314 => pixel <= "000000";
      when 7315 => pixel <= "000000";
      when 7316 => pixel <= "000000";
      when 7317 => pixel <= "000000";
      when 7318 => pixel <= "000000";
      when 7319 => pixel <= "001101";
      when 7320 => pixel <= "001101";
      when 7321 => pixel <= "000000";
      when 7322 => pixel <= "000000";
      when 7323 => pixel <= "000000";
      when 7324 => pixel <= "000000";
      when 7325 => pixel <= "001101";
      when 7326 => pixel <= "001101";
      when 7327 => pixel <= "000000";
      when 7328 => pixel <= "000000";
      when 7329 => pixel <= "000000";
      when 7330 => pixel <= "001101";
      when 7331 => pixel <= "001101";
      when 7332 => pixel <= "000000";
      when 7333 => pixel <= "000000";
      when 7334 => pixel <= "000000";
      when 7335 => pixel <= "000000";
      when 7336 => pixel <= "000000";
      when 7337 => pixel <= "000000";
      when 7338 => pixel <= "000000";
      when 7339 => pixel <= "000000";
      when 7340 => pixel <= "000000";
      when 7341 => pixel <= "000000";
      when 7342 => pixel <= "000000";
      when 7343 => pixel <= "000000";
      when 7344 => pixel <= "000000";
      when 7345 => pixel <= "000000";
      when 7346 => pixel <= "000000";
      when 7347 => pixel <= "000000";
      when 7348 => pixel <= "000000";
      when 7349 => pixel <= "000000";
      when 7350 => pixel <= "000000";
      when 7351 => pixel <= "000000";
      when 7352 => pixel <= "000000";
      when 7353 => pixel <= "000000";
      when 7354 => pixel <= "000000";
      when 7355 => pixel <= "000000";
      when 7356 => pixel <= "000000";
      when 7357 => pixel <= "000000";
      when 7358 => pixel <= "000000";
      when 7359 => pixel <= "000000";
      when 7360 => pixel <= "000000";
      when 7361 => pixel <= "000000";
      when 7362 => pixel <= "000000";
      when 7363 => pixel <= "000000";
      when 7364 => pixel <= "000000";
      when 7365 => pixel <= "000000";
      when 7366 => pixel <= "000000";
      when 7367 => pixel <= "000000";
      when 7368 => pixel <= "000000";
      when 7369 => pixel <= "000000";
      when 7370 => pixel <= "000000";
      when 7371 => pixel <= "000000";
      when 7372 => pixel <= "000000";
      when 7373 => pixel <= "000000";
      when 7374 => pixel <= "000000";
      when 7375 => pixel <= "000000";
      when 7376 => pixel <= "000000";
      when 7377 => pixel <= "000000";
      when 7378 => pixel <= "000000";
      when 7379 => pixel <= "000000";
      when 7380 => pixel <= "000000";
      when 7381 => pixel <= "000000";
      when 7382 => pixel <= "000000";
      when 7383 => pixel <= "000000";
      when 7384 => pixel <= "000000";
      when 7385 => pixel <= "000000";
      when 7386 => pixel <= "001101";
      when 7387 => pixel <= "001101";
      when 7388 => pixel <= "000000";
      when 7389 => pixel <= "000000";
      when 7390 => pixel <= "000000";
      when 7391 => pixel <= "000000";
      when 7392 => pixel <= "000000";
      when 7393 => pixel <= "000000";
      when 7394 => pixel <= "000000";
      when 7395 => pixel <= "001101";
      when 7396 => pixel <= "001101";
      when 7397 => pixel <= "000000";
      when 7398 => pixel <= "000000";
      when 7399 => pixel <= "001101";
      when 7400 => pixel <= "001101";
      when 7401 => pixel <= "000000";
      when 7402 => pixel <= "000000";
      when 7403 => pixel <= "000000";
      when 7404 => pixel <= "001101";
      when 7405 => pixel <= "001101";
      when 7406 => pixel <= "000000";
      when 7407 => pixel <= "000000";
      when 7408 => pixel <= "000000";
      when 7409 => pixel <= "001101";
      when 7410 => pixel <= "000000";
      when 7411 => pixel <= "000000";
      when 7412 => pixel <= "001101";
      when 7413 => pixel <= "001101";
      when 7414 => pixel <= "000000";
      when 7415 => pixel <= "000000";
      when 7416 => pixel <= "000000";
      when 7417 => pixel <= "001101";
      when 7418 => pixel <= "001101";
      when 7419 => pixel <= "000000";
      when 7420 => pixel <= "000000";
      when 7421 => pixel <= "001101";
      when 7422 => pixel <= "001101";
      when 7423 => pixel <= "000000";
      when 7424 => pixel <= "000000";
      when 7425 => pixel <= "000000";
      when 7426 => pixel <= "001101";
      when 7427 => pixel <= "001101";
      when 7428 => pixel <= "000000";
      when 7429 => pixel <= "000000";
      when 7430 => pixel <= "000000";
      when 7431 => pixel <= "000000";
      when 7432 => pixel <= "000000";
      when 7433 => pixel <= "000000";
      when 7434 => pixel <= "000000";
      when 7435 => pixel <= "000000";
      when 7436 => pixel <= "000000";
      when 7437 => pixel <= "000000";
      when 7438 => pixel <= "000000";
      when 7439 => pixel <= "000000";
      when 7440 => pixel <= "000000";
      when 7441 => pixel <= "000000";
      when 7442 => pixel <= "001101";
      when 7443 => pixel <= "001101";
      when 7444 => pixel <= "000000";
      when 7445 => pixel <= "000000";
      when 7446 => pixel <= "000000";
      when 7447 => pixel <= "000000";
      when 7448 => pixel <= "000000";
      when 7449 => pixel <= "001101";
      when 7450 => pixel <= "001101";
      when 7451 => pixel <= "000000";
      when 7452 => pixel <= "000000";
      when 7453 => pixel <= "000000";
      when 7454 => pixel <= "001101";
      when 7455 => pixel <= "001101";
      when 7456 => pixel <= "000000";
      when 7457 => pixel <= "000000";
      when 7458 => pixel <= "000000";
      when 7459 => pixel <= "000000";
      when 7460 => pixel <= "000000";
      when 7461 => pixel <= "000000";
      when 7462 => pixel <= "001101";
      when 7463 => pixel <= "001101";
      when 7464 => pixel <= "000000";
      when 7465 => pixel <= "000000";
      when 7466 => pixel <= "000000";
      when 7467 => pixel <= "000000";
      when 7468 => pixel <= "000000";
      when 7469 => pixel <= "000000";
      when 7470 => pixel <= "000000";
      when 7471 => pixel <= "000000";
      when 7472 => pixel <= "000000";
      when 7473 => pixel <= "000000";
      when 7474 => pixel <= "000000";
      when 7475 => pixel <= "000000";
      when 7476 => pixel <= "000000";
      when 7477 => pixel <= "000000";
      when 7478 => pixel <= "000000";
      when 7479 => pixel <= "001101";
      when 7480 => pixel <= "001101";
      when 7481 => pixel <= "000000";
      when 7482 => pixel <= "000000";
      when 7483 => pixel <= "000000";
      when 7484 => pixel <= "000000";
      when 7485 => pixel <= "001101";
      when 7486 => pixel <= "001101";
      when 7487 => pixel <= "000000";
      when 7488 => pixel <= "000000";
      when 7489 => pixel <= "000000";
      when 7490 => pixel <= "001101";
      when 7491 => pixel <= "001101";
      when 7492 => pixel <= "000000";
      when 7493 => pixel <= "000000";
      when 7494 => pixel <= "000000";
      when 7495 => pixel <= "000000";
      when 7496 => pixel <= "000000";
      when 7497 => pixel <= "000000";
      when 7498 => pixel <= "000000";
      when 7499 => pixel <= "000000";
      when 7500 => pixel <= "000000";
      when 7501 => pixel <= "000000";
      when 7502 => pixel <= "000000";
      when 7503 => pixel <= "000000";
      when 7504 => pixel <= "000000";
      when 7505 => pixel <= "000000";
      when 7506 => pixel <= "000000";
      when 7507 => pixel <= "000000";
      when 7508 => pixel <= "000000";
      when 7509 => pixel <= "000000";
      when 7510 => pixel <= "000000";
      when 7511 => pixel <= "000000";
      when 7512 => pixel <= "000000";
      when 7513 => pixel <= "000000";
      when 7514 => pixel <= "000000";
      when 7515 => pixel <= "000000";
      when 7516 => pixel <= "000000";
      when 7517 => pixel <= "000000";
      when 7518 => pixel <= "000000";
      when 7519 => pixel <= "000000";
      when 7520 => pixel <= "000000";
      when 7521 => pixel <= "000000";
      when 7522 => pixel <= "000000";
      when 7523 => pixel <= "000000";
      when 7524 => pixel <= "000000";
      when 7525 => pixel <= "000000";
      when 7526 => pixel <= "000000";
      when 7527 => pixel <= "000000";
      when 7528 => pixel <= "000000";
      when 7529 => pixel <= "000000";
      when 7530 => pixel <= "000000";
      when 7531 => pixel <= "000000";
      when 7532 => pixel <= "000000";
      when 7533 => pixel <= "000000";
      when 7534 => pixel <= "000000";
      when 7535 => pixel <= "000000";
      when 7536 => pixel <= "000000";
      when 7537 => pixel <= "000000";
      when 7538 => pixel <= "000000";
      when 7539 => pixel <= "000000";
      when 7540 => pixel <= "000000";
      when 7541 => pixel <= "000000";
      when 7542 => pixel <= "000000";
      when 7543 => pixel <= "000000";
      when 7544 => pixel <= "000000";
      when 7545 => pixel <= "000000";
      when 7546 => pixel <= "001101";
      when 7547 => pixel <= "001101";
      when 7548 => pixel <= "000000";
      when 7549 => pixel <= "000000";
      when 7550 => pixel <= "000000";
      when 7551 => pixel <= "000000";
      when 7552 => pixel <= "000000";
      when 7553 => pixel <= "000000";
      when 7554 => pixel <= "000000";
      when 7555 => pixel <= "001101";
      when 7556 => pixel <= "001101";
      when 7557 => pixel <= "000000";
      when 7558 => pixel <= "000000";
      when 7559 => pixel <= "001101";
      when 7560 => pixel <= "001101";
      when 7561 => pixel <= "000000";
      when 7562 => pixel <= "000000";
      when 7563 => pixel <= "000000";
      when 7564 => pixel <= "001101";
      when 7565 => pixel <= "001101";
      when 7566 => pixel <= "000000";
      when 7567 => pixel <= "000000";
      when 7568 => pixel <= "001101";
      when 7569 => pixel <= "001101";
      when 7570 => pixel <= "000000";
      when 7571 => pixel <= "000000";
      when 7572 => pixel <= "001101";
      when 7573 => pixel <= "001101";
      when 7574 => pixel <= "000000";
      when 7575 => pixel <= "000000";
      when 7576 => pixel <= "000000";
      when 7577 => pixel <= "001101";
      when 7578 => pixel <= "001101";
      when 7579 => pixel <= "000000";
      when 7580 => pixel <= "000000";
      when 7581 => pixel <= "001101";
      when 7582 => pixel <= "001101";
      when 7583 => pixel <= "000000";
      when 7584 => pixel <= "000000";
      when 7585 => pixel <= "000000";
      when 7586 => pixel <= "001101";
      when 7587 => pixel <= "001101";
      when 7588 => pixel <= "000000";
      when 7589 => pixel <= "000000";
      when 7590 => pixel <= "000000";
      when 7591 => pixel <= "000000";
      when 7592 => pixel <= "000000";
      when 7593 => pixel <= "000000";
      when 7594 => pixel <= "000000";
      when 7595 => pixel <= "000000";
      when 7596 => pixel <= "000000";
      when 7597 => pixel <= "000000";
      when 7598 => pixel <= "000000";
      when 7599 => pixel <= "000000";
      when 7600 => pixel <= "000000";
      when 7601 => pixel <= "000000";
      when 7602 => pixel <= "000000";
      when 7603 => pixel <= "001101";
      when 7604 => pixel <= "001101";
      when 7605 => pixel <= "000000";
      when 7606 => pixel <= "000000";
      when 7607 => pixel <= "000000";
      when 7608 => pixel <= "000000";
      when 7609 => pixel <= "001101";
      when 7610 => pixel <= "001101";
      when 7611 => pixel <= "000000";
      when 7612 => pixel <= "000000";
      when 7613 => pixel <= "000000";
      when 7614 => pixel <= "001101";
      when 7615 => pixel <= "001101";
      when 7616 => pixel <= "000000";
      when 7617 => pixel <= "000000";
      when 7618 => pixel <= "000000";
      when 7619 => pixel <= "000000";
      when 7620 => pixel <= "000000";
      when 7621 => pixel <= "001101";
      when 7622 => pixel <= "001101";
      when 7623 => pixel <= "000000";
      when 7624 => pixel <= "000000";
      when 7625 => pixel <= "000000";
      when 7626 => pixel <= "000000";
      when 7627 => pixel <= "000000";
      when 7628 => pixel <= "000000";
      when 7629 => pixel <= "000000";
      when 7630 => pixel <= "000000";
      when 7631 => pixel <= "000000";
      when 7632 => pixel <= "000000";
      when 7633 => pixel <= "000000";
      when 7634 => pixel <= "000000";
      when 7635 => pixel <= "000000";
      when 7636 => pixel <= "000000";
      when 7637 => pixel <= "000000";
      when 7638 => pixel <= "000000";
      when 7639 => pixel <= "001101";
      when 7640 => pixel <= "001101";
      when 7641 => pixel <= "000000";
      when 7642 => pixel <= "000000";
      when 7643 => pixel <= "000000";
      when 7644 => pixel <= "000000";
      when 7645 => pixel <= "001101";
      when 7646 => pixel <= "001101";
      when 7647 => pixel <= "000000";
      when 7648 => pixel <= "000000";
      when 7649 => pixel <= "000000";
      when 7650 => pixel <= "001101";
      when 7651 => pixel <= "001101";
      when 7652 => pixel <= "000000";
      when 7653 => pixel <= "000000";
      when 7654 => pixel <= "000000";
      when 7655 => pixel <= "000000";
      when 7656 => pixel <= "000000";
      when 7657 => pixel <= "000000";
      when 7658 => pixel <= "000000";
      when 7659 => pixel <= "000000";
      when 7660 => pixel <= "000000";
      when 7661 => pixel <= "000000";
      when 7662 => pixel <= "000000";
      when 7663 => pixel <= "000000";
      when 7664 => pixel <= "000000";
      when 7665 => pixel <= "000000";
      when 7666 => pixel <= "000000";
      when 7667 => pixel <= "000000";
      when 7668 => pixel <= "000000";
      when 7669 => pixel <= "000000";
      when 7670 => pixel <= "000000";
      when 7671 => pixel <= "000000";
      when 7672 => pixel <= "000000";
      when 7673 => pixel <= "000000";
      when 7674 => pixel <= "000000";
      when 7675 => pixel <= "000000";
      when 7676 => pixel <= "000000";
      when 7677 => pixel <= "000000";
      when 7678 => pixel <= "000000";
      when 7679 => pixel <= "000000";
      when 7680 => pixel <= "000000";
      when 7681 => pixel <= "000000";
      when 7682 => pixel <= "000000";
      when 7683 => pixel <= "000000";
      when 7684 => pixel <= "000000";
      when 7685 => pixel <= "000000";
      when 7686 => pixel <= "000000";
      when 7687 => pixel <= "000000";
      when 7688 => pixel <= "000000";
      when 7689 => pixel <= "000000";
      when 7690 => pixel <= "000000";
      when 7691 => pixel <= "000000";
      when 7692 => pixel <= "000000";
      when 7693 => pixel <= "000000";
      when 7694 => pixel <= "000000";
      when 7695 => pixel <= "000000";
      when 7696 => pixel <= "000000";
      when 7697 => pixel <= "000000";
      when 7698 => pixel <= "000000";
      when 7699 => pixel <= "000000";
      when 7700 => pixel <= "000000";
      when 7701 => pixel <= "000000";
      when 7702 => pixel <= "000000";
      when 7703 => pixel <= "000000";
      when 7704 => pixel <= "000000";
      when 7705 => pixel <= "001101";
      when 7706 => pixel <= "001101";
      when 7707 => pixel <= "001101";
      when 7708 => pixel <= "001101";
      when 7709 => pixel <= "000000";
      when 7710 => pixel <= "000000";
      when 7711 => pixel <= "000000";
      when 7712 => pixel <= "000000";
      when 7713 => pixel <= "000000";
      when 7714 => pixel <= "001101";
      when 7715 => pixel <= "001101";
      when 7716 => pixel <= "001101";
      when 7717 => pixel <= "000000";
      when 7718 => pixel <= "000000";
      when 7719 => pixel <= "001101";
      when 7720 => pixel <= "001101";
      when 7721 => pixel <= "000000";
      when 7722 => pixel <= "000000";
      when 7723 => pixel <= "001101";
      when 7724 => pixel <= "001101";
      when 7725 => pixel <= "001101";
      when 7726 => pixel <= "001101";
      when 7727 => pixel <= "001101";
      when 7728 => pixel <= "001101";
      when 7729 => pixel <= "001101";
      when 7730 => pixel <= "000000";
      when 7731 => pixel <= "000000";
      when 7732 => pixel <= "000000";
      when 7733 => pixel <= "001101";
      when 7734 => pixel <= "001101";
      when 7735 => pixel <= "001101";
      when 7736 => pixel <= "001101";
      when 7737 => pixel <= "001101";
      when 7738 => pixel <= "000000";
      when 7739 => pixel <= "000000";
      when 7740 => pixel <= "000000";
      when 7741 => pixel <= "000000";
      when 7742 => pixel <= "001101";
      when 7743 => pixel <= "001101";
      when 7744 => pixel <= "001101";
      when 7745 => pixel <= "001101";
      when 7746 => pixel <= "001101";
      when 7747 => pixel <= "000000";
      when 7748 => pixel <= "000000";
      when 7749 => pixel <= "000000";
      when 7750 => pixel <= "000000";
      when 7751 => pixel <= "000000";
      when 7752 => pixel <= "000000";
      when 7753 => pixel <= "000000";
      when 7754 => pixel <= "000000";
      when 7755 => pixel <= "000000";
      when 7756 => pixel <= "000000";
      when 7757 => pixel <= "000000";
      when 7758 => pixel <= "000000";
      when 7759 => pixel <= "000000";
      when 7760 => pixel <= "000000";
      when 7761 => pixel <= "000000";
      when 7762 => pixel <= "000000";
      when 7763 => pixel <= "000000";
      when 7764 => pixel <= "001101";
      when 7765 => pixel <= "001101";
      when 7766 => pixel <= "000000";
      when 7767 => pixel <= "000000";
      when 7768 => pixel <= "000000";
      when 7769 => pixel <= "001101";
      when 7770 => pixel <= "001101";
      when 7771 => pixel <= "000000";
      when 7772 => pixel <= "000000";
      when 7773 => pixel <= "000000";
      when 7774 => pixel <= "001101";
      when 7775 => pixel <= "001101";
      when 7776 => pixel <= "000000";
      when 7777 => pixel <= "000000";
      when 7778 => pixel <= "000000";
      when 7779 => pixel <= "000000";
      when 7780 => pixel <= "001101";
      when 7781 => pixel <= "001101";
      when 7782 => pixel <= "000000";
      when 7783 => pixel <= "000000";
      when 7784 => pixel <= "000000";
      when 7785 => pixel <= "000000";
      when 7786 => pixel <= "000000";
      when 7787 => pixel <= "000000";
      when 7788 => pixel <= "000000";
      when 7789 => pixel <= "000000";
      when 7790 => pixel <= "000000";
      when 7791 => pixel <= "000000";
      when 7792 => pixel <= "000000";
      when 7793 => pixel <= "000000";
      when 7794 => pixel <= "000000";
      when 7795 => pixel <= "000000";
      when 7796 => pixel <= "000000";
      when 7797 => pixel <= "000000";
      when 7798 => pixel <= "001101";
      when 7799 => pixel <= "001101";
      when 7800 => pixel <= "001101";
      when 7801 => pixel <= "001101";
      when 7802 => pixel <= "000000";
      when 7803 => pixel <= "000000";
      when 7804 => pixel <= "000000";
      when 7805 => pixel <= "000000";
      when 7806 => pixel <= "001101";
      when 7807 => pixel <= "001101";
      when 7808 => pixel <= "001101";
      when 7809 => pixel <= "001101";
      when 7810 => pixel <= "001101";
      when 7811 => pixel <= "000000";
      when 7812 => pixel <= "000000";
      when 7813 => pixel <= "000000";
      when 7814 => pixel <= "000000";
      when 7815 => pixel <= "000000";
      when 7816 => pixel <= "000000";
      when 7817 => pixel <= "000000";
      when 7818 => pixel <= "000000";
      when 7819 => pixel <= "000000";
      when 7820 => pixel <= "000000";
      when 7821 => pixel <= "000000";
      when 7822 => pixel <= "000000";
      when 7823 => pixel <= "000000";
      when 7824 => pixel <= "000000";
      when 7825 => pixel <= "000000";
      when 7826 => pixel <= "000000";
      when 7827 => pixel <= "000000";
      when 7828 => pixel <= "000000";
      when 7829 => pixel <= "000000";
      when 7830 => pixel <= "000000";
      when 7831 => pixel <= "000000";
      when 7832 => pixel <= "000000";
      when 7833 => pixel <= "000000";
      when 7834 => pixel <= "000000";
      when 7835 => pixel <= "000000";
      when 7836 => pixel <= "000000";
      when 7837 => pixel <= "000000";
      when 7838 => pixel <= "000000";
      when 7839 => pixel <= "000000";
      when 7840 => pixel <= "000000";
      when 7841 => pixel <= "000000";
      when 7842 => pixel <= "000000";
      when 7843 => pixel <= "000000";
      when 7844 => pixel <= "000000";
      when 7845 => pixel <= "000000";
      when 7846 => pixel <= "000000";
      when 7847 => pixel <= "000000";
      when 7848 => pixel <= "000000";
      when 7849 => pixel <= "000000";
      when 7850 => pixel <= "000000";
      when 7851 => pixel <= "000000";
      when 7852 => pixel <= "000000";
      when 7853 => pixel <= "000000";
      when 7854 => pixel <= "000000";
      when 7855 => pixel <= "000000";
      when 7856 => pixel <= "000000";
      when 7857 => pixel <= "000000";
      when 7858 => pixel <= "000000";
      when 7859 => pixel <= "000000";
      when 7860 => pixel <= "000000";
      when 7861 => pixel <= "000000";
      when 7862 => pixel <= "000000";
      when 7863 => pixel <= "000000";
      when 7864 => pixel <= "000000";
      when 7865 => pixel <= "000000";
      when 7866 => pixel <= "000000";
      when 7867 => pixel <= "000000";
      when 7868 => pixel <= "000000";
      when 7869 => pixel <= "000000";
      when 7870 => pixel <= "000000";
      when 7871 => pixel <= "000000";
      when 7872 => pixel <= "000000";
      when 7873 => pixel <= "000000";
      when 7874 => pixel <= "000000";
      when 7875 => pixel <= "000000";
      when 7876 => pixel <= "000000";
      when 7877 => pixel <= "000000";
      when 7878 => pixel <= "000000";
      when 7879 => pixel <= "000000";
      when 7880 => pixel <= "000000";
      when 7881 => pixel <= "000000";
      when 7882 => pixel <= "000000";
      when 7883 => pixel <= "000000";
      when 7884 => pixel <= "000000";
      when 7885 => pixel <= "000000";
      when 7886 => pixel <= "000000";
      when 7887 => pixel <= "000000";
      when 7888 => pixel <= "000000";
      when 7889 => pixel <= "000000";
      when 7890 => pixel <= "000000";
      when 7891 => pixel <= "000000";
      when 7892 => pixel <= "000000";
      when 7893 => pixel <= "000000";
      when 7894 => pixel <= "000000";
      when 7895 => pixel <= "000000";
      when 7896 => pixel <= "000000";
      when 7897 => pixel <= "000000";
      when 7898 => pixel <= "000000";
      when 7899 => pixel <= "000000";
      when 7900 => pixel <= "000000";
      when 7901 => pixel <= "000000";
      when 7902 => pixel <= "000000";
      when 7903 => pixel <= "000000";
      when 7904 => pixel <= "000000";
      when 7905 => pixel <= "000000";
      when 7906 => pixel <= "000000";
      when 7907 => pixel <= "000000";
      when 7908 => pixel <= "000000";
      when 7909 => pixel <= "000000";
      when 7910 => pixel <= "000000";
      when 7911 => pixel <= "000000";
      when 7912 => pixel <= "000000";
      when 7913 => pixel <= "000000";
      when 7914 => pixel <= "000000";
      when 7915 => pixel <= "000000";
      when 7916 => pixel <= "000000";
      when 7917 => pixel <= "000000";
      when 7918 => pixel <= "000000";
      when 7919 => pixel <= "000000";
      when 7920 => pixel <= "000000";
      when 7921 => pixel <= "000000";
      when 7922 => pixel <= "000000";
      when 7923 => pixel <= "000000";
      when 7924 => pixel <= "000000";
      when 7925 => pixel <= "000000";
      when 7926 => pixel <= "000000";
      when 7927 => pixel <= "000000";
      when 7928 => pixel <= "000000";
      when 7929 => pixel <= "000000";
      when 7930 => pixel <= "000000";
      when 7931 => pixel <= "000000";
      when 7932 => pixel <= "000000";
      when 7933 => pixel <= "000000";
      when 7934 => pixel <= "000000";
      when 7935 => pixel <= "000000";
      when 7936 => pixel <= "000000";
      when 7937 => pixel <= "000000";
      when 7938 => pixel <= "000000";
      when 7939 => pixel <= "000000";
      when 7940 => pixel <= "000000";
      when 7941 => pixel <= "000000";
      when 7942 => pixel <= "000000";
      when 7943 => pixel <= "000000";
      when 7944 => pixel <= "000000";
      when 7945 => pixel <= "000000";
      when 7946 => pixel <= "000000";
      when 7947 => pixel <= "000000";
      when 7948 => pixel <= "000000";
      when 7949 => pixel <= "000000";
      when 7950 => pixel <= "000000";
      when 7951 => pixel <= "000000";
      when 7952 => pixel <= "000000";
      when 7953 => pixel <= "000000";
      when 7954 => pixel <= "000000";
      when 7955 => pixel <= "000000";
      when 7956 => pixel <= "000000";
      when 7957 => pixel <= "000000";
      when 7958 => pixel <= "000000";
      when 7959 => pixel <= "000000";
      when 7960 => pixel <= "000000";
      when 7961 => pixel <= "000000";
      when 7962 => pixel <= "000000";
      when 7963 => pixel <= "000000";
      when 7964 => pixel <= "000000";
      when 7965 => pixel <= "000000";
      when 7966 => pixel <= "000000";
      when 7967 => pixel <= "000000";
      when 7968 => pixel <= "000000";
      when 7969 => pixel <= "000000";
      when 7970 => pixel <= "000000";
      when 7971 => pixel <= "000000";
      when 7972 => pixel <= "000000";
      when 7973 => pixel <= "000000";
      when 7974 => pixel <= "000000";
      when 7975 => pixel <= "000000";
      when 7976 => pixel <= "000000";
      when 7977 => pixel <= "000000";
      when 7978 => pixel <= "000000";
      when 7979 => pixel <= "000000";
      when 7980 => pixel <= "000000";
      when 7981 => pixel <= "000000";
      when 7982 => pixel <= "000000";
      when 7983 => pixel <= "000000";
      when 7984 => pixel <= "000000";
      when 7985 => pixel <= "000000";
      when 7986 => pixel <= "000000";
      when 7987 => pixel <= "000000";
      when 7988 => pixel <= "000000";
      when 7989 => pixel <= "000000";
      when 7990 => pixel <= "000000";
      when 7991 => pixel <= "000000";
      when 7992 => pixel <= "000000";
      when 7993 => pixel <= "000000";
      when 7994 => pixel <= "000000";
      when 7995 => pixel <= "000000";
      when 7996 => pixel <= "000000";
      when 7997 => pixel <= "000000";
      when 7998 => pixel <= "000000";
      when 7999 => pixel <= "000000";
      when 8000 => pixel <= "000000";
      when 8001 => pixel <= "000000";
      when 8002 => pixel <= "000000";
      when 8003 => pixel <= "000000";
      when 8004 => pixel <= "000000";
      when 8005 => pixel <= "000000";
      when 8006 => pixel <= "000000";
      when 8007 => pixel <= "000000";
      when 8008 => pixel <= "000000";
      when 8009 => pixel <= "000000";
      when 8010 => pixel <= "000000";
      when 8011 => pixel <= "000000";
      when 8012 => pixel <= "000000";
      when 8013 => pixel <= "000000";
      when 8014 => pixel <= "000000";
      when 8015 => pixel <= "000000";
      when 8016 => pixel <= "000000";
      when 8017 => pixel <= "000000";
      when 8018 => pixel <= "000000";
      when 8019 => pixel <= "000000";
      when 8020 => pixel <= "000000";
      when 8021 => pixel <= "000000";
      when 8022 => pixel <= "000000";
      when 8023 => pixel <= "000000";
      when 8024 => pixel <= "000000";
      when 8025 => pixel <= "000000";
      when 8026 => pixel <= "000000";
      when 8027 => pixel <= "000000";
      when 8028 => pixel <= "000000";
      when 8029 => pixel <= "000000";
      when 8030 => pixel <= "000000";
      when 8031 => pixel <= "000000";
      when 8032 => pixel <= "000000";
      when 8033 => pixel <= "000000";
      when 8034 => pixel <= "000000";
      when 8035 => pixel <= "000000";
      when 8036 => pixel <= "000000";
      when 8037 => pixel <= "000000";
      when 8038 => pixel <= "000000";
      when 8039 => pixel <= "000000";
      when 8040 => pixel <= "000000";
      when 8041 => pixel <= "000000";
      when 8042 => pixel <= "000000";
      when 8043 => pixel <= "000000";
      when 8044 => pixel <= "000000";
      when 8045 => pixel <= "000000";
      when 8046 => pixel <= "000000";
      when 8047 => pixel <= "000000";
      when 8048 => pixel <= "000000";
      when 8049 => pixel <= "000000";
      when 8050 => pixel <= "000000";
      when 8051 => pixel <= "000000";
      when 8052 => pixel <= "000000";
      when 8053 => pixel <= "000000";
      when 8054 => pixel <= "000000";
      when 8055 => pixel <= "000000";
      when 8056 => pixel <= "000000";
      when 8057 => pixel <= "000000";
      when 8058 => pixel <= "000000";
      when 8059 => pixel <= "000000";
      when 8060 => pixel <= "000000";
      when 8061 => pixel <= "000000";
      when 8062 => pixel <= "000000";
      when 8063 => pixel <= "000000";
      when 8064 => pixel <= "000000";
      when 8065 => pixel <= "000000";
      when 8066 => pixel <= "000000";
      when 8067 => pixel <= "000000";
      when 8068 => pixel <= "000000";
      when 8069 => pixel <= "000000";
      when 8070 => pixel <= "000000";
      when 8071 => pixel <= "000000";
      when 8072 => pixel <= "000000";
      when 8073 => pixel <= "000000";
      when 8074 => pixel <= "000000";
      when 8075 => pixel <= "000000";
      when 8076 => pixel <= "000000";
      when 8077 => pixel <= "000000";
      when 8078 => pixel <= "000000";
      when 8079 => pixel <= "000000";
      when 8080 => pixel <= "000000";
      when 8081 => pixel <= "000000";
      when 8082 => pixel <= "000000";
      when 8083 => pixel <= "000000";
      when 8084 => pixel <= "000000";
      when 8085 => pixel <= "000000";
      when 8086 => pixel <= "000000";
      when 8087 => pixel <= "000000";
      when 8088 => pixel <= "000000";
      when 8089 => pixel <= "000000";
      when 8090 => pixel <= "000000";
      when 8091 => pixel <= "000000";
      when 8092 => pixel <= "000000";
      when 8093 => pixel <= "000000";
      when 8094 => pixel <= "000000";
      when 8095 => pixel <= "000000";
      when 8096 => pixel <= "000000";
      when 8097 => pixel <= "000000";
      when 8098 => pixel <= "000000";
      when 8099 => pixel <= "000000";
      when 8100 => pixel <= "000000";
      when 8101 => pixel <= "000000";
      when 8102 => pixel <= "000000";
      when 8103 => pixel <= "000000";
      when 8104 => pixel <= "000000";
      when 8105 => pixel <= "000000";
      when 8106 => pixel <= "000000";
      when 8107 => pixel <= "000000";
      when 8108 => pixel <= "000000";
      when 8109 => pixel <= "000000";
      when 8110 => pixel <= "000000";
      when 8111 => pixel <= "000000";
      when 8112 => pixel <= "000000";
      when 8113 => pixel <= "000000";
      when 8114 => pixel <= "000000";
      when 8115 => pixel <= "000000";
      when 8116 => pixel <= "000000";
      when 8117 => pixel <= "000000";
      when 8118 => pixel <= "000000";
      when 8119 => pixel <= "000000";
      when 8120 => pixel <= "000000";
      when 8121 => pixel <= "000000";
      when 8122 => pixel <= "000000";
      when 8123 => pixel <= "000000";
      when 8124 => pixel <= "000000";
      when 8125 => pixel <= "000000";
      when 8126 => pixel <= "000000";
      when 8127 => pixel <= "000000";
      when 8128 => pixel <= "000000";
      when 8129 => pixel <= "000000";
      when 8130 => pixel <= "000000";
      when 8131 => pixel <= "000000";
      when 8132 => pixel <= "000000";
      when 8133 => pixel <= "000000";
      when 8134 => pixel <= "000000";
      when 8135 => pixel <= "000000";
      when 8136 => pixel <= "000000";
      when 8137 => pixel <= "000000";
      when 8138 => pixel <= "000000";
      when 8139 => pixel <= "000000";
      when 8140 => pixel <= "000000";
      when 8141 => pixel <= "000000";
      when 8142 => pixel <= "000000";
      when 8143 => pixel <= "000000";
      when 8144 => pixel <= "000000";
      when 8145 => pixel <= "000000";
      when 8146 => pixel <= "000000";
      when 8147 => pixel <= "000000";
      when 8148 => pixel <= "000000";
      when 8149 => pixel <= "000000";
      when 8150 => pixel <= "000000";
      when 8151 => pixel <= "000000";
      when 8152 => pixel <= "000000";
      when 8153 => pixel <= "000000";
      when 8154 => pixel <= "000000";
      when 8155 => pixel <= "000000";
      when 8156 => pixel <= "000000";
      when 8157 => pixel <= "000000";
      when 8158 => pixel <= "000000";
      when 8159 => pixel <= "000000";
      when 8160 => pixel <= "000000";
      when 8161 => pixel <= "000000";
      when 8162 => pixel <= "000000";
      when 8163 => pixel <= "000000";
      when 8164 => pixel <= "000000";
      when 8165 => pixel <= "000000";
      when 8166 => pixel <= "000000";
      when 8167 => pixel <= "000000";
      when 8168 => pixel <= "000000";
      when 8169 => pixel <= "000000";
      when 8170 => pixel <= "000000";
      when 8171 => pixel <= "000000";
      when 8172 => pixel <= "000000";
      when 8173 => pixel <= "000000";
      when 8174 => pixel <= "000000";
      when 8175 => pixel <= "000000";
      when 8176 => pixel <= "000000";
      when 8177 => pixel <= "000000";
      when 8178 => pixel <= "000000";
      when 8179 => pixel <= "000000";
      when 8180 => pixel <= "000000";
      when 8181 => pixel <= "000000";
      when 8182 => pixel <= "000000";
      when 8183 => pixel <= "000000";
      when 8184 => pixel <= "000000";
      when 8185 => pixel <= "000000";
      when 8186 => pixel <= "000000";
      when 8187 => pixel <= "000000";
      when 8188 => pixel <= "000000";
      when 8189 => pixel <= "000000";
      when 8190 => pixel <= "000000";
      when 8191 => pixel <= "000000";
      when 8192 => pixel <= "000000";
      when 8193 => pixel <= "000000";
      when 8194 => pixel <= "000000";
      when 8195 => pixel <= "000000";
      when 8196 => pixel <= "000000";
      when 8197 => pixel <= "000000";
      when 8198 => pixel <= "000000";
      when 8199 => pixel <= "000000";
      when 8200 => pixel <= "000000";
      when 8201 => pixel <= "000000";
      when 8202 => pixel <= "000000";
      when 8203 => pixel <= "000000";
      when 8204 => pixel <= "000000";
      when 8205 => pixel <= "000000";
      when 8206 => pixel <= "000000";
      when 8207 => pixel <= "000000";
      when 8208 => pixel <= "000000";
      when 8209 => pixel <= "000000";
      when 8210 => pixel <= "000000";
      when 8211 => pixel <= "000000";
      when 8212 => pixel <= "000000";
      when 8213 => pixel <= "000000";
      when 8214 => pixel <= "000000";
      when 8215 => pixel <= "000000";
      when 8216 => pixel <= "000000";
      when 8217 => pixel <= "000000";
      when 8218 => pixel <= "000000";
      when 8219 => pixel <= "000000";
      when 8220 => pixel <= "000000";
      when 8221 => pixel <= "000000";
      when 8222 => pixel <= "000000";
      when 8223 => pixel <= "000000";
      when 8224 => pixel <= "000000";
      when 8225 => pixel <= "000000";
      when 8226 => pixel <= "000000";
      when 8227 => pixel <= "000000";
      when 8228 => pixel <= "000000";
      when 8229 => pixel <= "000000";
      when 8230 => pixel <= "000000";
      when 8231 => pixel <= "000000";
      when 8232 => pixel <= "000000";
      when 8233 => pixel <= "000000";
      when 8234 => pixel <= "000000";
      when 8235 => pixel <= "000000";
      when 8236 => pixel <= "000000";
      when 8237 => pixel <= "000000";
      when 8238 => pixel <= "000000";
      when 8239 => pixel <= "000000";
      when 8240 => pixel <= "000000";
      when 8241 => pixel <= "000000";
      when 8242 => pixel <= "000000";
      when 8243 => pixel <= "000000";
      when 8244 => pixel <= "000000";
      when 8245 => pixel <= "000000";
      when 8246 => pixel <= "000000";
      when 8247 => pixel <= "000000";
      when 8248 => pixel <= "000000";
      when 8249 => pixel <= "000000";
      when 8250 => pixel <= "000000";
      when 8251 => pixel <= "000000";
      when 8252 => pixel <= "000000";
      when 8253 => pixel <= "000000";
      when 8254 => pixel <= "000000";
      when 8255 => pixel <= "000000";
      when 8256 => pixel <= "000000";
      when 8257 => pixel <= "000000";
      when 8258 => pixel <= "000000";
      when 8259 => pixel <= "000000";
      when 8260 => pixel <= "000000";
      when 8261 => pixel <= "000000";
      when 8262 => pixel <= "000000";
      when 8263 => pixel <= "000000";
      when 8264 => pixel <= "000000";
      when 8265 => pixel <= "000000";
      when 8266 => pixel <= "000000";
      when 8267 => pixel <= "000000";
      when 8268 => pixel <= "000000";
      when 8269 => pixel <= "000000";
      when 8270 => pixel <= "000000";
      when 8271 => pixel <= "000000";
      when 8272 => pixel <= "000000";
      when 8273 => pixel <= "000000";
      when 8274 => pixel <= "000000";
      when 8275 => pixel <= "000000";
      when 8276 => pixel <= "000000";
      when 8277 => pixel <= "000000";
      when 8278 => pixel <= "000000";
      when 8279 => pixel <= "000000";
      when 8280 => pixel <= "000000";
      when 8281 => pixel <= "000000";
      when 8282 => pixel <= "000000";
      when 8283 => pixel <= "000000";
      when 8284 => pixel <= "000000";
      when 8285 => pixel <= "000000";
      when 8286 => pixel <= "000000";
      when 8287 => pixel <= "000000";
      when 8288 => pixel <= "000000";
      when 8289 => pixel <= "000000";
      when 8290 => pixel <= "000000";
      when 8291 => pixel <= "000000";
      when 8292 => pixel <= "000000";
      when 8293 => pixel <= "000000";
      when 8294 => pixel <= "000000";
      when 8295 => pixel <= "000000";
      when 8296 => pixel <= "000000";
      when 8297 => pixel <= "000000";
      when 8298 => pixel <= "000000";
      when 8299 => pixel <= "000000";
      when 8300 => pixel <= "000000";
      when 8301 => pixel <= "000000";
      when 8302 => pixel <= "000000";
      when 8303 => pixel <= "000000";
      when 8304 => pixel <= "000000";
      when 8305 => pixel <= "000000";
      when 8306 => pixel <= "000000";
      when 8307 => pixel <= "000000";
      when 8308 => pixel <= "000000";
      when 8309 => pixel <= "000000";
      when 8310 => pixel <= "000000";
      when 8311 => pixel <= "000000";
      when 8312 => pixel <= "000000";
      when 8313 => pixel <= "000000";
      when 8314 => pixel <= "000000";
      when 8315 => pixel <= "000000";
      when 8316 => pixel <= "000000";
      when 8317 => pixel <= "000000";
      when 8318 => pixel <= "000000";
      when 8319 => pixel <= "000000";
      when 8320 => pixel <= "000000";
      when 8321 => pixel <= "000000";
      when 8322 => pixel <= "000000";
      when 8323 => pixel <= "000000";
      when 8324 => pixel <= "000000";
      when 8325 => pixel <= "000000";
      when 8326 => pixel <= "000000";
      when 8327 => pixel <= "000000";
      when 8328 => pixel <= "000000";
      when 8329 => pixel <= "000000";
      when 8330 => pixel <= "000000";
      when 8331 => pixel <= "000000";
      when 8332 => pixel <= "000000";
      when 8333 => pixel <= "000000";
      when 8334 => pixel <= "000000";
      when 8335 => pixel <= "000000";
      when 8336 => pixel <= "000000";
      when 8337 => pixel <= "000000";
      when 8338 => pixel <= "000000";
      when 8339 => pixel <= "000000";
      when 8340 => pixel <= "000000";
      when 8341 => pixel <= "000000";
      when 8342 => pixel <= "000000";
      when 8343 => pixel <= "000000";
      when 8344 => pixel <= "000000";
      when 8345 => pixel <= "000000";
      when 8346 => pixel <= "000000";
      when 8347 => pixel <= "000000";
      when 8348 => pixel <= "000000";
      when 8349 => pixel <= "000000";
      when 8350 => pixel <= "000000";
      when 8351 => pixel <= "000000";
      when 8352 => pixel <= "000000";
      when 8353 => pixel <= "000000";
      when 8354 => pixel <= "000000";
      when 8355 => pixel <= "000000";
      when 8356 => pixel <= "000000";
      when 8357 => pixel <= "000000";
      when 8358 => pixel <= "000000";
      when 8359 => pixel <= "000000";
      when 8360 => pixel <= "000000";
      when 8361 => pixel <= "000000";
      when 8362 => pixel <= "000000";
      when 8363 => pixel <= "000000";
      when 8364 => pixel <= "000000";
      when 8365 => pixel <= "000000";
      when 8366 => pixel <= "000000";
      when 8367 => pixel <= "000000";
      when 8368 => pixel <= "000000";
      when 8369 => pixel <= "000000";
      when 8370 => pixel <= "000000";
      when 8371 => pixel <= "000000";
      when 8372 => pixel <= "000000";
      when 8373 => pixel <= "000000";
      when 8374 => pixel <= "000000";
      when 8375 => pixel <= "000000";
      when 8376 => pixel <= "000000";
      when 8377 => pixel <= "000000";
      when 8378 => pixel <= "000000";
      when 8379 => pixel <= "000000";
      when 8380 => pixel <= "000000";
      when 8381 => pixel <= "000000";
      when 8382 => pixel <= "000000";
      when 8383 => pixel <= "000000";
      when 8384 => pixel <= "000000";
      when 8385 => pixel <= "000000";
      when 8386 => pixel <= "000000";
      when 8387 => pixel <= "000000";
      when 8388 => pixel <= "000000";
      when 8389 => pixel <= "000000";
      when 8390 => pixel <= "000000";
      when 8391 => pixel <= "000000";
      when 8392 => pixel <= "000000";
      when 8393 => pixel <= "000000";
      when 8394 => pixel <= "000000";
      when 8395 => pixel <= "000000";
      when 8396 => pixel <= "000000";
      when 8397 => pixel <= "000000";
      when 8398 => pixel <= "000000";
      when 8399 => pixel <= "000000";
      when 8400 => pixel <= "000000";
      when 8401 => pixel <= "000000";
      when 8402 => pixel <= "000000";
      when 8403 => pixel <= "000000";
      when 8404 => pixel <= "000000";
      when 8405 => pixel <= "000000";
      when 8406 => pixel <= "000000";
      when 8407 => pixel <= "000000";
      when 8408 => pixel <= "000000";
      when 8409 => pixel <= "000000";
      when 8410 => pixel <= "000000";
      when 8411 => pixel <= "000000";
      when 8412 => pixel <= "000000";
      when 8413 => pixel <= "000000";
      when 8414 => pixel <= "000000";
      when 8415 => pixel <= "000000";
      when 8416 => pixel <= "000000";
      when 8417 => pixel <= "000000";
      when 8418 => pixel <= "000000";
      when 8419 => pixel <= "000000";
      when 8420 => pixel <= "000000";
      when 8421 => pixel <= "000000";
      when 8422 => pixel <= "000000";
      when 8423 => pixel <= "000000";
      when 8424 => pixel <= "000000";
      when 8425 => pixel <= "000000";
      when 8426 => pixel <= "000000";
      when 8427 => pixel <= "000000";
      when 8428 => pixel <= "000000";
      when 8429 => pixel <= "000000";
      when 8430 => pixel <= "000000";
      when 8431 => pixel <= "000000";
      when 8432 => pixel <= "000000";
      when 8433 => pixel <= "000000";
      when 8434 => pixel <= "000000";
      when 8435 => pixel <= "000000";
      when 8436 => pixel <= "000000";
      when 8437 => pixel <= "000000";
      when 8438 => pixel <= "000000";
      when 8439 => pixel <= "000000";
      when 8440 => pixel <= "000000";
      when 8441 => pixel <= "000000";
      when 8442 => pixel <= "000000";
      when 8443 => pixel <= "000000";
      when 8444 => pixel <= "000000";
      when 8445 => pixel <= "000000";
      when 8446 => pixel <= "000000";
      when 8447 => pixel <= "000000";
      when 8448 => pixel <= "000000";
      when 8449 => pixel <= "000000";
      when 8450 => pixel <= "000000";
      when 8451 => pixel <= "000000";
      when 8452 => pixel <= "000000";
      when 8453 => pixel <= "000000";
      when 8454 => pixel <= "000000";
      when 8455 => pixel <= "000000";
      when 8456 => pixel <= "000000";
      when 8457 => pixel <= "000000";
      when 8458 => pixel <= "000000";
      when 8459 => pixel <= "000000";
      when 8460 => pixel <= "000000";
      when 8461 => pixel <= "000000";
      when 8462 => pixel <= "000000";
      when 8463 => pixel <= "000000";
      when 8464 => pixel <= "000000";
      when 8465 => pixel <= "000000";
      when 8466 => pixel <= "000000";
      when 8467 => pixel <= "000000";
      when 8468 => pixel <= "000000";
      when 8469 => pixel <= "000000";
      when 8470 => pixel <= "000000";
      when 8471 => pixel <= "000000";
      when 8472 => pixel <= "000000";
      when 8473 => pixel <= "000000";
      when 8474 => pixel <= "000000";
      when 8475 => pixel <= "000000";
      when 8476 => pixel <= "000000";
      when 8477 => pixel <= "000000";
      when 8478 => pixel <= "000000";
      when 8479 => pixel <= "000000";
      when 8480 => pixel <= "000000";
      when 8481 => pixel <= "000000";
      when 8482 => pixel <= "000000";
      when 8483 => pixel <= "000000";
      when 8484 => pixel <= "000000";
      when 8485 => pixel <= "000000";
      when 8486 => pixel <= "000000";
      when 8487 => pixel <= "000000";
      when 8488 => pixel <= "000000";
      when 8489 => pixel <= "000000";
      when 8490 => pixel <= "000000";
      when 8491 => pixel <= "000000";
      when 8492 => pixel <= "000000";
      when 8493 => pixel <= "000000";
      when 8494 => pixel <= "000000";
      when 8495 => pixel <= "000000";
      when 8496 => pixel <= "000000";
      when 8497 => pixel <= "000000";
      when 8498 => pixel <= "000000";
      when 8499 => pixel <= "000000";
      when 8500 => pixel <= "000000";
      when 8501 => pixel <= "000000";
      when 8502 => pixel <= "000000";
      when 8503 => pixel <= "000000";
      when 8504 => pixel <= "000000";
      when 8505 => pixel <= "000000";
      when 8506 => pixel <= "000000";
      when 8507 => pixel <= "000000";
      when 8508 => pixel <= "000000";
      when 8509 => pixel <= "000000";
      when 8510 => pixel <= "000000";
      when 8511 => pixel <= "000000";
      when 8512 => pixel <= "000000";
      when 8513 => pixel <= "000000";
      when 8514 => pixel <= "000000";
      when 8515 => pixel <= "000000";
      when 8516 => pixel <= "000000";
      when 8517 => pixel <= "000000";
      when 8518 => pixel <= "000000";
      when 8519 => pixel <= "000000";
      when 8520 => pixel <= "000000";
      when 8521 => pixel <= "000000";
      when 8522 => pixel <= "000000";
      when 8523 => pixel <= "000000";
      when 8524 => pixel <= "000000";
      when 8525 => pixel <= "000000";
      when 8526 => pixel <= "000000";
      when 8527 => pixel <= "000000";
      when 8528 => pixel <= "000000";
      when 8529 => pixel <= "000000";
      when 8530 => pixel <= "000000";
      when 8531 => pixel <= "000000";
      when 8532 => pixel <= "000000";
      when 8533 => pixel <= "000000";
      when 8534 => pixel <= "000000";
      when 8535 => pixel <= "000000";
      when 8536 => pixel <= "000000";
      when 8537 => pixel <= "000000";
      when 8538 => pixel <= "000000";
      when 8539 => pixel <= "000000";
      when 8540 => pixel <= "000000";
      when 8541 => pixel <= "000000";
      when 8542 => pixel <= "000000";
      when 8543 => pixel <= "000000";
      when 8544 => pixel <= "000000";
      when 8545 => pixel <= "000000";
      when 8546 => pixel <= "000000";
      when 8547 => pixel <= "000000";
      when 8548 => pixel <= "000000";
      when 8549 => pixel <= "000000";
      when 8550 => pixel <= "000000";
      when 8551 => pixel <= "000000";
      when 8552 => pixel <= "000000";
      when 8553 => pixel <= "000000";
      when 8554 => pixel <= "000000";
      when 8555 => pixel <= "000000";
      when 8556 => pixel <= "000000";
      when 8557 => pixel <= "000000";
      when 8558 => pixel <= "000000";
      when 8559 => pixel <= "000000";
      when 8560 => pixel <= "000000";
      when 8561 => pixel <= "000000";
      when 8562 => pixel <= "000000";
      when 8563 => pixel <= "000000";
      when 8564 => pixel <= "000000";
      when 8565 => pixel <= "000000";
      when 8566 => pixel <= "000000";
      when 8567 => pixel <= "000000";
      when 8568 => pixel <= "000000";
      when 8569 => pixel <= "000000";
      when 8570 => pixel <= "000000";
      when 8571 => pixel <= "000000";
      when 8572 => pixel <= "000000";
      when 8573 => pixel <= "000000";
      when 8574 => pixel <= "000000";
      when 8575 => pixel <= "000000";
      when 8576 => pixel <= "000000";
      when 8577 => pixel <= "000000";
      when 8578 => pixel <= "000000";
      when 8579 => pixel <= "000000";
      when 8580 => pixel <= "000000";
      when 8581 => pixel <= "000000";
      when 8582 => pixel <= "000000";
      when 8583 => pixel <= "000000";
      when 8584 => pixel <= "000000";
      when 8585 => pixel <= "000000";
      when 8586 => pixel <= "000000";
      when 8587 => pixel <= "000000";
      when 8588 => pixel <= "000000";
      when 8589 => pixel <= "000000";
      when 8590 => pixel <= "000000";
      when 8591 => pixel <= "000000";
      when 8592 => pixel <= "000000";
      when 8593 => pixel <= "000000";
      when 8594 => pixel <= "000000";
      when 8595 => pixel <= "000000";
      when 8596 => pixel <= "000000";
      when 8597 => pixel <= "000000";
      when 8598 => pixel <= "000000";
      when 8599 => pixel <= "000000";
      when 8600 => pixel <= "000000";
      when 8601 => pixel <= "000000";
      when 8602 => pixel <= "000000";
      when 8603 => pixel <= "000000";
      when 8604 => pixel <= "000000";
      when 8605 => pixel <= "000000";
      when 8606 => pixel <= "000000";
      when 8607 => pixel <= "000000";
      when 8608 => pixel <= "000000";
      when 8609 => pixel <= "000000";
      when 8610 => pixel <= "000000";
      when 8611 => pixel <= "000000";
      when 8612 => pixel <= "000000";
      when 8613 => pixel <= "000000";
      when 8614 => pixel <= "000000";
      when 8615 => pixel <= "000000";
      when 8616 => pixel <= "000000";
      when 8617 => pixel <= "000000";
      when 8618 => pixel <= "000000";
      when 8619 => pixel <= "000000";
      when 8620 => pixel <= "000000";
      when 8621 => pixel <= "000000";
      when 8622 => pixel <= "000000";
      when 8623 => pixel <= "000000";
      when 8624 => pixel <= "000000";
      when 8625 => pixel <= "000000";
      when 8626 => pixel <= "000000";
      when 8627 => pixel <= "000000";
      when 8628 => pixel <= "000000";
      when 8629 => pixel <= "000000";
      when 8630 => pixel <= "000000";
      when 8631 => pixel <= "000000";
      when 8632 => pixel <= "000000";
      when 8633 => pixel <= "000000";
      when 8634 => pixel <= "000000";
      when 8635 => pixel <= "000000";
      when 8636 => pixel <= "000000";
      when 8637 => pixel <= "000000";
      when 8638 => pixel <= "000000";
      when 8639 => pixel <= "000000";
      when 8640 => pixel <= "000000";
      when 8641 => pixel <= "000000";
      when 8642 => pixel <= "000000";
      when 8643 => pixel <= "000000";
      when 8644 => pixel <= "000000";
      when 8645 => pixel <= "000000";
      when 8646 => pixel <= "000000";
      when 8647 => pixel <= "000000";
      when 8648 => pixel <= "000000";
      when 8649 => pixel <= "000000";
      when 8650 => pixel <= "000000";
      when 8651 => pixel <= "000000";
      when 8652 => pixel <= "000000";
      when 8653 => pixel <= "000000";
      when 8654 => pixel <= "000000";
      when 8655 => pixel <= "000000";
      when 8656 => pixel <= "000000";
      when 8657 => pixel <= "000000";
      when 8658 => pixel <= "000000";
      when 8659 => pixel <= "000000";
      when 8660 => pixel <= "000000";
      when 8661 => pixel <= "000000";
      when 8662 => pixel <= "000000";
      when 8663 => pixel <= "000000";
      when 8664 => pixel <= "000000";
      when 8665 => pixel <= "000000";
      when 8666 => pixel <= "000000";
      when 8667 => pixel <= "000000";
      when 8668 => pixel <= "000000";
      when 8669 => pixel <= "000000";
      when 8670 => pixel <= "000000";
      when 8671 => pixel <= "000000";
      when 8672 => pixel <= "000000";
      when 8673 => pixel <= "000000";
      when 8674 => pixel <= "000000";
      when 8675 => pixel <= "000000";
      when 8676 => pixel <= "000000";
      when 8677 => pixel <= "000000";
      when 8678 => pixel <= "000000";
      when 8679 => pixel <= "000000";
      when 8680 => pixel <= "000000";
      when 8681 => pixel <= "000000";
      when 8682 => pixel <= "000000";
      when 8683 => pixel <= "000000";
      when 8684 => pixel <= "000000";
      when 8685 => pixel <= "000000";
      when 8686 => pixel <= "000000";
      when 8687 => pixel <= "000000";
      when 8688 => pixel <= "000000";
      when 8689 => pixel <= "000000";
      when 8690 => pixel <= "000000";
      when 8691 => pixel <= "000000";
      when 8692 => pixel <= "000000";
      when 8693 => pixel <= "000000";
      when 8694 => pixel <= "000000";
      when 8695 => pixel <= "000000";
      when 8696 => pixel <= "000000";
      when 8697 => pixel <= "000000";
      when 8698 => pixel <= "000000";
      when 8699 => pixel <= "000000";
      when 8700 => pixel <= "000000";
      when 8701 => pixel <= "000000";
      when 8702 => pixel <= "000000";
      when 8703 => pixel <= "000000";
      when 8704 => pixel <= "000000";
      when 8705 => pixel <= "000000";
      when 8706 => pixel <= "000000";
      when 8707 => pixel <= "000000";
      when 8708 => pixel <= "000000";
      when 8709 => pixel <= "000000";
      when 8710 => pixel <= "000000";
      when 8711 => pixel <= "000000";
      when 8712 => pixel <= "000000";
      when 8713 => pixel <= "000000";
      when 8714 => pixel <= "000000";
      when 8715 => pixel <= "000000";
      when 8716 => pixel <= "000000";
      when 8717 => pixel <= "000000";
      when 8718 => pixel <= "000000";
      when 8719 => pixel <= "000000";
      when 8720 => pixel <= "000000";
      when 8721 => pixel <= "000000";
      when 8722 => pixel <= "000000";
      when 8723 => pixel <= "000000";
      when 8724 => pixel <= "000000";
      when 8725 => pixel <= "000000";
      when 8726 => pixel <= "000000";
      when 8727 => pixel <= "000000";
      when 8728 => pixel <= "000000";
      when 8729 => pixel <= "000000";
      when 8730 => pixel <= "000000";
      when 8731 => pixel <= "000000";
      when 8732 => pixel <= "000000";
      when 8733 => pixel <= "000000";
      when 8734 => pixel <= "000000";
      when 8735 => pixel <= "000000";
      when 8736 => pixel <= "000000";
      when 8737 => pixel <= "000000";
      when 8738 => pixel <= "000000";
      when 8739 => pixel <= "000000";
      when 8740 => pixel <= "000000";
      when 8741 => pixel <= "000000";
      when 8742 => pixel <= "000000";
      when 8743 => pixel <= "000000";
      when 8744 => pixel <= "000000";
      when 8745 => pixel <= "000000";
      when 8746 => pixel <= "000000";
      when 8747 => pixel <= "000000";
      when 8748 => pixel <= "000000";
      when 8749 => pixel <= "000000";
      when 8750 => pixel <= "000000";
      when 8751 => pixel <= "000000";
      when 8752 => pixel <= "000000";
      when 8753 => pixel <= "000000";
      when 8754 => pixel <= "000000";
      when 8755 => pixel <= "000000";
      when 8756 => pixel <= "000000";
      when 8757 => pixel <= "000000";
      when 8758 => pixel <= "000000";
      when 8759 => pixel <= "000000";
      when 8760 => pixel <= "000000";
      when 8761 => pixel <= "000000";
      when 8762 => pixel <= "000000";
      when 8763 => pixel <= "000000";
      when 8764 => pixel <= "000000";
      when 8765 => pixel <= "000000";
      when 8766 => pixel <= "000000";
      when 8767 => pixel <= "000000";
      when 8768 => pixel <= "000000";
      when 8769 => pixel <= "000000";
      when 8770 => pixel <= "000000";
      when 8771 => pixel <= "000000";
      when 8772 => pixel <= "000000";
      when 8773 => pixel <= "000000";
      when 8774 => pixel <= "000000";
      when 8775 => pixel <= "000000";
      when 8776 => pixel <= "000000";
      when 8777 => pixel <= "000000";
      when 8778 => pixel <= "000000";
      when 8779 => pixel <= "000000";
      when 8780 => pixel <= "000000";
      when 8781 => pixel <= "000000";
      when 8782 => pixel <= "000000";
      when 8783 => pixel <= "000000";
      when 8784 => pixel <= "000000";
      when 8785 => pixel <= "000000";
      when 8786 => pixel <= "000000";
      when 8787 => pixel <= "000000";
      when 8788 => pixel <= "000000";
      when 8789 => pixel <= "000000";
      when 8790 => pixel <= "000000";
      when 8791 => pixel <= "000000";
      when 8792 => pixel <= "000000";
      when 8793 => pixel <= "000000";
      when 8794 => pixel <= "000000";
      when 8795 => pixel <= "000000";
      when 8796 => pixel <= "000000";
      when 8797 => pixel <= "000000";
      when 8798 => pixel <= "000000";
      when 8799 => pixel <= "000000";
      when 8800 => pixel <= "000000";
      when 8801 => pixel <= "000000";
      when 8802 => pixel <= "000000";
      when 8803 => pixel <= "000000";
      when 8804 => pixel <= "000000";
      when 8805 => pixel <= "000000";
      when 8806 => pixel <= "000000";
      when 8807 => pixel <= "000000";
      when 8808 => pixel <= "000000";
      when 8809 => pixel <= "000000";
      when 8810 => pixel <= "000000";
      when 8811 => pixel <= "000000";
      when 8812 => pixel <= "000000";
      when 8813 => pixel <= "000000";
      when 8814 => pixel <= "000000";
      when 8815 => pixel <= "000000";
      when 8816 => pixel <= "000000";
      when 8817 => pixel <= "000000";
      when 8818 => pixel <= "000000";
      when 8819 => pixel <= "000000";
      when 8820 => pixel <= "000000";
      when 8821 => pixel <= "000000";
      when 8822 => pixel <= "000000";
      when 8823 => pixel <= "000000";
      when 8824 => pixel <= "000000";
      when 8825 => pixel <= "000000";
      when 8826 => pixel <= "000000";
      when 8827 => pixel <= "000000";
      when 8828 => pixel <= "000000";
      when 8829 => pixel <= "000000";
      when 8830 => pixel <= "000000";
      when 8831 => pixel <= "000000";
      when 8832 => pixel <= "000000";
      when 8833 => pixel <= "000000";
      when 8834 => pixel <= "001101";
      when 8835 => pixel <= "001101";
      when 8836 => pixel <= "001101";
      when 8837 => pixel <= "001101";
      when 8838 => pixel <= "001101";
      when 8839 => pixel <= "001101";
      when 8840 => pixel <= "000000";
      when 8841 => pixel <= "000000";
      when 8842 => pixel <= "000000";
      when 8843 => pixel <= "001101";
      when 8844 => pixel <= "001101";
      when 8845 => pixel <= "001101";
      when 8846 => pixel <= "001101";
      when 8847 => pixel <= "000000";
      when 8848 => pixel <= "000000";
      when 8849 => pixel <= "000000";
      when 8850 => pixel <= "000000";
      when 8851 => pixel <= "000000";
      when 8852 => pixel <= "000000";
      when 8853 => pixel <= "000000";
      when 8854 => pixel <= "000000";
      when 8855 => pixel <= "001101";
      when 8856 => pixel <= "000000";
      when 8857 => pixel <= "000000";
      when 8858 => pixel <= "000000";
      when 8859 => pixel <= "000000";
      when 8860 => pixel <= "000000";
      when 8861 => pixel <= "000000";
      when 8862 => pixel <= "001101";
      when 8863 => pixel <= "001101";
      when 8864 => pixel <= "000000";
      when 8865 => pixel <= "000000";
      when 8866 => pixel <= "001101";
      when 8867 => pixel <= "001101";
      when 8868 => pixel <= "000000";
      when 8869 => pixel <= "000000";
      when 8870 => pixel <= "000000";
      when 8871 => pixel <= "000000";
      when 8872 => pixel <= "000000";
      when 8873 => pixel <= "000000";
      when 8874 => pixel <= "000000";
      when 8875 => pixel <= "000000";
      when 8876 => pixel <= "000000";
      when 8877 => pixel <= "000000";
      when 8878 => pixel <= "000000";
      when 8879 => pixel <= "000000";
      when 8880 => pixel <= "000000";
      when 8881 => pixel <= "000000";
      when 8882 => pixel <= "000000";
      when 8883 => pixel <= "001101";
      when 8884 => pixel <= "000000";
      when 8885 => pixel <= "000000";
      when 8886 => pixel <= "000000";
      when 8887 => pixel <= "000000";
      when 8888 => pixel <= "000000";
      when 8889 => pixel <= "000000";
      when 8890 => pixel <= "000000";
      when 8891 => pixel <= "001101";
      when 8892 => pixel <= "001101";
      when 8893 => pixel <= "001101";
      when 8894 => pixel <= "001101";
      when 8895 => pixel <= "000000";
      when 8896 => pixel <= "000000";
      when 8897 => pixel <= "000000";
      when 8898 => pixel <= "000000";
      when 8899 => pixel <= "000000";
      when 8900 => pixel <= "000000";
      when 8901 => pixel <= "001101";
      when 8902 => pixel <= "000000";
      when 8903 => pixel <= "000000";
      when 8904 => pixel <= "000000";
      when 8905 => pixel <= "000000";
      when 8906 => pixel <= "000000";
      when 8907 => pixel <= "000000";
      when 8908 => pixel <= "000000";
      when 8909 => pixel <= "001101";
      when 8910 => pixel <= "001101";
      when 8911 => pixel <= "001101";
      when 8912 => pixel <= "001101";
      when 8913 => pixel <= "000000";
      when 8914 => pixel <= "000000";
      when 8915 => pixel <= "000000";
      when 8916 => pixel <= "001101";
      when 8917 => pixel <= "001101";
      when 8918 => pixel <= "000000";
      when 8919 => pixel <= "000000";
      when 8920 => pixel <= "000000";
      when 8921 => pixel <= "001101";
      when 8922 => pixel <= "001101";
      when 8923 => pixel <= "000000";
      when 8924 => pixel <= "000000";
      when 8925 => pixel <= "000000";
      when 8926 => pixel <= "000000";
      when 8927 => pixel <= "000000";
      when 8928 => pixel <= "000000";
      when 8929 => pixel <= "000000";
      when 8930 => pixel <= "000000";
      when 8931 => pixel <= "000000";
      when 8932 => pixel <= "000000";
      when 8933 => pixel <= "000000";
      when 8934 => pixel <= "000000";
      when 8935 => pixel <= "000000";
      when 8936 => pixel <= "000000";
      when 8937 => pixel <= "000000";
      when 8938 => pixel <= "000000";
      when 8939 => pixel <= "000000";
      when 8940 => pixel <= "000000";
      when 8941 => pixel <= "000000";
      when 8942 => pixel <= "000000";
      when 8943 => pixel <= "000000";
      when 8944 => pixel <= "000000";
      when 8945 => pixel <= "000000";
      when 8946 => pixel <= "000000";
      when 8947 => pixel <= "000000";
      when 8948 => pixel <= "000000";
      when 8949 => pixel <= "000000";
      when 8950 => pixel <= "000000";
      when 8951 => pixel <= "000000";
      when 8952 => pixel <= "000000";
      when 8953 => pixel <= "000000";
      when 8954 => pixel <= "000000";
      when 8955 => pixel <= "000000";
      when 8956 => pixel <= "000000";
      when 8957 => pixel <= "000000";
      when 8958 => pixel <= "000000";
      when 8959 => pixel <= "000000";
      when 8960 => pixel <= "000000";
      when 8961 => pixel <= "000000";
      when 8962 => pixel <= "000000";
      when 8963 => pixel <= "000000";
      when 8964 => pixel <= "000000";
      when 8965 => pixel <= "000000";
      when 8966 => pixel <= "000000";
      when 8967 => pixel <= "000000";
      when 8968 => pixel <= "000000";
      when 8969 => pixel <= "000000";
      when 8970 => pixel <= "000000";
      when 8971 => pixel <= "000000";
      when 8972 => pixel <= "000000";
      when 8973 => pixel <= "000000";
      when 8974 => pixel <= "000000";
      when 8975 => pixel <= "000000";
      when 8976 => pixel <= "000000";
      when 8977 => pixel <= "000000";
      when 8978 => pixel <= "000000";
      when 8979 => pixel <= "000000";
      when 8980 => pixel <= "000000";
      when 8981 => pixel <= "000000";
      when 8982 => pixel <= "000000";
      when 8983 => pixel <= "000000";
      when 8984 => pixel <= "000000";
      when 8985 => pixel <= "000000";
      when 8986 => pixel <= "000000";
      when 8987 => pixel <= "000000";
      when 8988 => pixel <= "000000";
      when 8989 => pixel <= "000000";
      when 8990 => pixel <= "000000";
      when 8991 => pixel <= "000000";
      when 8992 => pixel <= "000000";
      when 8993 => pixel <= "000000";
      when 8994 => pixel <= "000000";
      when 8995 => pixel <= "001101";
      when 8996 => pixel <= "001101";
      when 8997 => pixel <= "000000";
      when 8998 => pixel <= "000000";
      when 8999 => pixel <= "001101";
      when 9000 => pixel <= "001101";
      when 9001 => pixel <= "000000";
      when 9002 => pixel <= "000000";
      when 9003 => pixel <= "000000";
      when 9004 => pixel <= "001101";
      when 9005 => pixel <= "001101";
      when 9006 => pixel <= "000000";
      when 9007 => pixel <= "000000";
      when 9008 => pixel <= "000000";
      when 9009 => pixel <= "000000";
      when 9010 => pixel <= "000000";
      when 9011 => pixel <= "000000";
      when 9012 => pixel <= "000000";
      when 9013 => pixel <= "000000";
      when 9014 => pixel <= "001101";
      when 9015 => pixel <= "001101";
      when 9016 => pixel <= "001101";
      when 9017 => pixel <= "000000";
      when 9018 => pixel <= "000000";
      when 9019 => pixel <= "000000";
      when 9020 => pixel <= "000000";
      when 9021 => pixel <= "000000";
      when 9022 => pixel <= "001101";
      when 9023 => pixel <= "001101";
      when 9024 => pixel <= "000000";
      when 9025 => pixel <= "000000";
      when 9026 => pixel <= "001101";
      when 9027 => pixel <= "001101";
      when 9028 => pixel <= "000000";
      when 9029 => pixel <= "000000";
      when 9030 => pixel <= "000000";
      when 9031 => pixel <= "000000";
      when 9032 => pixel <= "000000";
      when 9033 => pixel <= "000000";
      when 9034 => pixel <= "000000";
      when 9035 => pixel <= "000000";
      when 9036 => pixel <= "000000";
      when 9037 => pixel <= "000000";
      when 9038 => pixel <= "000000";
      when 9039 => pixel <= "000000";
      when 9040 => pixel <= "000000";
      when 9041 => pixel <= "000000";
      when 9042 => pixel <= "001101";
      when 9043 => pixel <= "001101";
      when 9044 => pixel <= "001101";
      when 9045 => pixel <= "000000";
      when 9046 => pixel <= "000000";
      when 9047 => pixel <= "000000";
      when 9048 => pixel <= "000000";
      when 9049 => pixel <= "000000";
      when 9050 => pixel <= "001101";
      when 9051 => pixel <= "001101";
      when 9052 => pixel <= "000000";
      when 9053 => pixel <= "000000";
      when 9054 => pixel <= "001101";
      when 9055 => pixel <= "001101";
      when 9056 => pixel <= "000000";
      when 9057 => pixel <= "000000";
      when 9058 => pixel <= "000000";
      when 9059 => pixel <= "000000";
      when 9060 => pixel <= "001101";
      when 9061 => pixel <= "001101";
      when 9062 => pixel <= "001101";
      when 9063 => pixel <= "000000";
      when 9064 => pixel <= "000000";
      when 9065 => pixel <= "000000";
      when 9066 => pixel <= "000000";
      when 9067 => pixel <= "000000";
      when 9068 => pixel <= "000000";
      when 9069 => pixel <= "000000";
      when 9070 => pixel <= "001101";
      when 9071 => pixel <= "001101";
      when 9072 => pixel <= "000000";
      when 9073 => pixel <= "000000";
      when 9074 => pixel <= "000000";
      when 9075 => pixel <= "000000";
      when 9076 => pixel <= "001101";
      when 9077 => pixel <= "001101";
      when 9078 => pixel <= "001101";
      when 9079 => pixel <= "000000";
      when 9080 => pixel <= "000000";
      when 9081 => pixel <= "001101";
      when 9082 => pixel <= "001101";
      when 9083 => pixel <= "000000";
      when 9084 => pixel <= "000000";
      when 9085 => pixel <= "000000";
      when 9086 => pixel <= "000000";
      when 9087 => pixel <= "000000";
      when 9088 => pixel <= "000000";
      when 9089 => pixel <= "000000";
      when 9090 => pixel <= "000000";
      when 9091 => pixel <= "000000";
      when 9092 => pixel <= "000000";
      when 9093 => pixel <= "000000";
      when 9094 => pixel <= "000000";
      when 9095 => pixel <= "000000";
      when 9096 => pixel <= "000000";
      when 9097 => pixel <= "000000";
      when 9098 => pixel <= "000000";
      when 9099 => pixel <= "000000";
      when 9100 => pixel <= "000000";
      when 9101 => pixel <= "000000";
      when 9102 => pixel <= "000000";
      when 9103 => pixel <= "000000";
      when 9104 => pixel <= "000000";
      when 9105 => pixel <= "000000";
      when 9106 => pixel <= "000000";
      when 9107 => pixel <= "000000";
      when 9108 => pixel <= "000000";
      when 9109 => pixel <= "000000";
      when 9110 => pixel <= "000000";
      when 9111 => pixel <= "000000";
      when 9112 => pixel <= "000000";
      when 9113 => pixel <= "000000";
      when 9114 => pixel <= "000000";
      when 9115 => pixel <= "000000";
      when 9116 => pixel <= "000000";
      when 9117 => pixel <= "000000";
      when 9118 => pixel <= "000000";
      when 9119 => pixel <= "000000";
      when 9120 => pixel <= "000000";
      when 9121 => pixel <= "000000";
      when 9122 => pixel <= "000000";
      when 9123 => pixel <= "000000";
      when 9124 => pixel <= "000000";
      when 9125 => pixel <= "000000";
      when 9126 => pixel <= "000000";
      when 9127 => pixel <= "000000";
      when 9128 => pixel <= "000000";
      when 9129 => pixel <= "000000";
      when 9130 => pixel <= "000000";
      when 9131 => pixel <= "000000";
      when 9132 => pixel <= "000000";
      when 9133 => pixel <= "000000";
      when 9134 => pixel <= "000000";
      when 9135 => pixel <= "000000";
      when 9136 => pixel <= "000000";
      when 9137 => pixel <= "000000";
      when 9138 => pixel <= "000000";
      when 9139 => pixel <= "000000";
      when 9140 => pixel <= "000000";
      when 9141 => pixel <= "000000";
      when 9142 => pixel <= "000000";
      when 9143 => pixel <= "000000";
      when 9144 => pixel <= "000000";
      when 9145 => pixel <= "000000";
      when 9146 => pixel <= "000000";
      when 9147 => pixel <= "000000";
      when 9148 => pixel <= "000000";
      when 9149 => pixel <= "000000";
      when 9150 => pixel <= "000000";
      when 9151 => pixel <= "000000";
      when 9152 => pixel <= "000000";
      when 9153 => pixel <= "000000";
      when 9154 => pixel <= "000000";
      when 9155 => pixel <= "001101";
      when 9156 => pixel <= "001101";
      when 9157 => pixel <= "000000";
      when 9158 => pixel <= "000000";
      when 9159 => pixel <= "001101";
      when 9160 => pixel <= "001101";
      when 9161 => pixel <= "000000";
      when 9162 => pixel <= "000000";
      when 9163 => pixel <= "000000";
      when 9164 => pixel <= "001101";
      when 9165 => pixel <= "001101";
      when 9166 => pixel <= "000000";
      when 9167 => pixel <= "000000";
      when 9168 => pixel <= "000000";
      when 9169 => pixel <= "000000";
      when 9170 => pixel <= "000000";
      when 9171 => pixel <= "000000";
      when 9172 => pixel <= "000000";
      when 9173 => pixel <= "001101";
      when 9174 => pixel <= "001101";
      when 9175 => pixel <= "000000";
      when 9176 => pixel <= "001101";
      when 9177 => pixel <= "001101";
      when 9178 => pixel <= "000000";
      when 9179 => pixel <= "000000";
      when 9180 => pixel <= "000000";
      when 9181 => pixel <= "000000";
      when 9182 => pixel <= "001101";
      when 9183 => pixel <= "001101";
      when 9184 => pixel <= "000000";
      when 9185 => pixel <= "000000";
      when 9186 => pixel <= "001101";
      when 9187 => pixel <= "001101";
      when 9188 => pixel <= "000000";
      when 9189 => pixel <= "000000";
      when 9190 => pixel <= "000000";
      when 9191 => pixel <= "000000";
      when 9192 => pixel <= "000000";
      when 9193 => pixel <= "000000";
      when 9194 => pixel <= "000000";
      when 9195 => pixel <= "000000";
      when 9196 => pixel <= "000000";
      when 9197 => pixel <= "000000";
      when 9198 => pixel <= "000000";
      when 9199 => pixel <= "000000";
      when 9200 => pixel <= "000000";
      when 9201 => pixel <= "001101";
      when 9202 => pixel <= "001101";
      when 9203 => pixel <= "000000";
      when 9204 => pixel <= "001101";
      when 9205 => pixel <= "001101";
      when 9206 => pixel <= "000000";
      when 9207 => pixel <= "000000";
      when 9208 => pixel <= "000000";
      when 9209 => pixel <= "001101";
      when 9210 => pixel <= "001101";
      when 9211 => pixel <= "000000";
      when 9212 => pixel <= "000000";
      when 9213 => pixel <= "000000";
      when 9214 => pixel <= "000000";
      when 9215 => pixel <= "001101";
      when 9216 => pixel <= "000000";
      when 9217 => pixel <= "000000";
      when 9218 => pixel <= "000000";
      when 9219 => pixel <= "001101";
      when 9220 => pixel <= "001101";
      when 9221 => pixel <= "000000";
      when 9222 => pixel <= "001101";
      when 9223 => pixel <= "001101";
      when 9224 => pixel <= "000000";
      when 9225 => pixel <= "000000";
      when 9226 => pixel <= "000000";
      when 9227 => pixel <= "000000";
      when 9228 => pixel <= "000000";
      when 9229 => pixel <= "000000";
      when 9230 => pixel <= "001101";
      when 9231 => pixel <= "001101";
      when 9232 => pixel <= "000000";
      when 9233 => pixel <= "000000";
      when 9234 => pixel <= "000000";
      when 9235 => pixel <= "000000";
      when 9236 => pixel <= "001101";
      when 9237 => pixel <= "001101";
      when 9238 => pixel <= "001101";
      when 9239 => pixel <= "001101";
      when 9240 => pixel <= "000000";
      when 9241 => pixel <= "001101";
      when 9242 => pixel <= "001101";
      when 9243 => pixel <= "000000";
      when 9244 => pixel <= "000000";
      when 9245 => pixel <= "000000";
      when 9246 => pixel <= "000000";
      when 9247 => pixel <= "000000";
      when 9248 => pixel <= "000000";
      when 9249 => pixel <= "000000";
      when 9250 => pixel <= "000000";
      when 9251 => pixel <= "000000";
      when 9252 => pixel <= "000000";
      when 9253 => pixel <= "000000";
      when 9254 => pixel <= "000000";
      when 9255 => pixel <= "000000";
      when 9256 => pixel <= "000000";
      when 9257 => pixel <= "000000";
      when 9258 => pixel <= "000000";
      when 9259 => pixel <= "000000";
      when 9260 => pixel <= "000000";
      when 9261 => pixel <= "000000";
      when 9262 => pixel <= "000000";
      when 9263 => pixel <= "000000";
      when 9264 => pixel <= "000000";
      when 9265 => pixel <= "000000";
      when 9266 => pixel <= "000000";
      when 9267 => pixel <= "000000";
      when 9268 => pixel <= "000000";
      when 9269 => pixel <= "000000";
      when 9270 => pixel <= "000000";
      when 9271 => pixel <= "000000";
      when 9272 => pixel <= "000000";
      when 9273 => pixel <= "000000";
      when 9274 => pixel <= "000000";
      when 9275 => pixel <= "000000";
      when 9276 => pixel <= "000000";
      when 9277 => pixel <= "000000";
      when 9278 => pixel <= "000000";
      when 9279 => pixel <= "000000";
      when 9280 => pixel <= "000000";
      when 9281 => pixel <= "000000";
      when 9282 => pixel <= "000000";
      when 9283 => pixel <= "000000";
      when 9284 => pixel <= "000000";
      when 9285 => pixel <= "000000";
      when 9286 => pixel <= "000000";
      when 9287 => pixel <= "000000";
      when 9288 => pixel <= "000000";
      when 9289 => pixel <= "000000";
      when 9290 => pixel <= "000000";
      when 9291 => pixel <= "000000";
      when 9292 => pixel <= "000000";
      when 9293 => pixel <= "000000";
      when 9294 => pixel <= "000000";
      when 9295 => pixel <= "000000";
      when 9296 => pixel <= "000000";
      when 9297 => pixel <= "000000";
      when 9298 => pixel <= "000000";
      when 9299 => pixel <= "000000";
      when 9300 => pixel <= "000000";
      when 9301 => pixel <= "000000";
      when 9302 => pixel <= "000000";
      when 9303 => pixel <= "000000";
      when 9304 => pixel <= "000000";
      when 9305 => pixel <= "000000";
      when 9306 => pixel <= "000000";
      when 9307 => pixel <= "000000";
      when 9308 => pixel <= "000000";
      when 9309 => pixel <= "000000";
      when 9310 => pixel <= "000000";
      when 9311 => pixel <= "000000";
      when 9312 => pixel <= "000000";
      when 9313 => pixel <= "000000";
      when 9314 => pixel <= "000000";
      when 9315 => pixel <= "001101";
      when 9316 => pixel <= "001101";
      when 9317 => pixel <= "000000";
      when 9318 => pixel <= "000000";
      when 9319 => pixel <= "001101";
      when 9320 => pixel <= "001101";
      when 9321 => pixel <= "000000";
      when 9322 => pixel <= "000000";
      when 9323 => pixel <= "000000";
      when 9324 => pixel <= "001101";
      when 9325 => pixel <= "001101";
      when 9326 => pixel <= "000000";
      when 9327 => pixel <= "000000";
      when 9328 => pixel <= "000000";
      when 9329 => pixel <= "000000";
      when 9330 => pixel <= "000000";
      when 9331 => pixel <= "000000";
      when 9332 => pixel <= "001101";
      when 9333 => pixel <= "001101";
      when 9334 => pixel <= "000000";
      when 9335 => pixel <= "000000";
      when 9336 => pixel <= "000000";
      when 9337 => pixel <= "001101";
      when 9338 => pixel <= "001101";
      when 9339 => pixel <= "000000";
      when 9340 => pixel <= "000000";
      when 9341 => pixel <= "000000";
      when 9342 => pixel <= "001101";
      when 9343 => pixel <= "001101";
      when 9344 => pixel <= "000000";
      when 9345 => pixel <= "000000";
      when 9346 => pixel <= "001101";
      when 9347 => pixel <= "001101";
      when 9348 => pixel <= "000000";
      when 9349 => pixel <= "000000";
      when 9350 => pixel <= "000000";
      when 9351 => pixel <= "000000";
      when 9352 => pixel <= "000000";
      when 9353 => pixel <= "000000";
      when 9354 => pixel <= "000000";
      when 9355 => pixel <= "000000";
      when 9356 => pixel <= "000000";
      when 9357 => pixel <= "000000";
      when 9358 => pixel <= "000000";
      when 9359 => pixel <= "001101";
      when 9360 => pixel <= "001101";
      when 9361 => pixel <= "001101";
      when 9362 => pixel <= "000000";
      when 9363 => pixel <= "000000";
      when 9364 => pixel <= "000000";
      when 9365 => pixel <= "001101";
      when 9366 => pixel <= "001101";
      when 9367 => pixel <= "000000";
      when 9368 => pixel <= "000000";
      when 9369 => pixel <= "001101";
      when 9370 => pixel <= "001101";
      when 9371 => pixel <= "000000";
      when 9372 => pixel <= "000000";
      when 9373 => pixel <= "000000";
      when 9374 => pixel <= "000000";
      when 9375 => pixel <= "000000";
      when 9376 => pixel <= "000000";
      when 9377 => pixel <= "000000";
      when 9378 => pixel <= "001101";
      when 9379 => pixel <= "001101";
      when 9380 => pixel <= "000000";
      when 9381 => pixel <= "000000";
      when 9382 => pixel <= "000000";
      when 9383 => pixel <= "001101";
      when 9384 => pixel <= "001101";
      when 9385 => pixel <= "000000";
      when 9386 => pixel <= "000000";
      when 9387 => pixel <= "000000";
      when 9388 => pixel <= "000000";
      when 9389 => pixel <= "000000";
      when 9390 => pixel <= "001101";
      when 9391 => pixel <= "001101";
      when 9392 => pixel <= "000000";
      when 9393 => pixel <= "000000";
      when 9394 => pixel <= "000000";
      when 9395 => pixel <= "000000";
      when 9396 => pixel <= "001101";
      when 9397 => pixel <= "001101";
      when 9398 => pixel <= "001101";
      when 9399 => pixel <= "001101";
      when 9400 => pixel <= "001101";
      when 9401 => pixel <= "001101";
      when 9402 => pixel <= "001101";
      when 9403 => pixel <= "000000";
      when 9404 => pixel <= "000000";
      when 9405 => pixel <= "000000";
      when 9406 => pixel <= "000000";
      when 9407 => pixel <= "000000";
      when 9408 => pixel <= "000000";
      when 9409 => pixel <= "000000";
      when 9410 => pixel <= "000000";
      when 9411 => pixel <= "000000";
      when 9412 => pixel <= "000000";
      when 9413 => pixel <= "000000";
      when 9414 => pixel <= "000000";
      when 9415 => pixel <= "000000";
      when 9416 => pixel <= "000000";
      when 9417 => pixel <= "000000";
      when 9418 => pixel <= "000000";
      when 9419 => pixel <= "000000";
      when 9420 => pixel <= "000000";
      when 9421 => pixel <= "000000";
      when 9422 => pixel <= "000000";
      when 9423 => pixel <= "000000";
      when 9424 => pixel <= "000000";
      when 9425 => pixel <= "000000";
      when 9426 => pixel <= "000000";
      when 9427 => pixel <= "000000";
      when 9428 => pixel <= "000000";
      when 9429 => pixel <= "000000";
      when 9430 => pixel <= "000000";
      when 9431 => pixel <= "000000";
      when 9432 => pixel <= "000000";
      when 9433 => pixel <= "000000";
      when 9434 => pixel <= "000000";
      when 9435 => pixel <= "000000";
      when 9436 => pixel <= "000000";
      when 9437 => pixel <= "000000";
      when 9438 => pixel <= "000000";
      when 9439 => pixel <= "000000";
      when 9440 => pixel <= "000000";
      when 9441 => pixel <= "000000";
      when 9442 => pixel <= "000000";
      when 9443 => pixel <= "000000";
      when 9444 => pixel <= "000000";
      when 9445 => pixel <= "000000";
      when 9446 => pixel <= "000000";
      when 9447 => pixel <= "000000";
      when 9448 => pixel <= "000000";
      when 9449 => pixel <= "000000";
      when 9450 => pixel <= "000000";
      when 9451 => pixel <= "000000";
      when 9452 => pixel <= "000000";
      when 9453 => pixel <= "000000";
      when 9454 => pixel <= "000000";
      when 9455 => pixel <= "000000";
      when 9456 => pixel <= "000000";
      when 9457 => pixel <= "000000";
      when 9458 => pixel <= "000000";
      when 9459 => pixel <= "000000";
      when 9460 => pixel <= "000000";
      when 9461 => pixel <= "000000";
      when 9462 => pixel <= "000000";
      when 9463 => pixel <= "000000";
      when 9464 => pixel <= "000000";
      when 9465 => pixel <= "000000";
      when 9466 => pixel <= "000000";
      when 9467 => pixel <= "000000";
      when 9468 => pixel <= "000000";
      when 9469 => pixel <= "000000";
      when 9470 => pixel <= "000000";
      when 9471 => pixel <= "000000";
      when 9472 => pixel <= "000000";
      when 9473 => pixel <= "000000";
      when 9474 => pixel <= "000000";
      when 9475 => pixel <= "001101";
      when 9476 => pixel <= "001101";
      when 9477 => pixel <= "001101";
      when 9478 => pixel <= "001101";
      when 9479 => pixel <= "001101";
      when 9480 => pixel <= "000000";
      when 9481 => pixel <= "000000";
      when 9482 => pixel <= "000000";
      when 9483 => pixel <= "000000";
      when 9484 => pixel <= "001101";
      when 9485 => pixel <= "001101";
      when 9486 => pixel <= "000000";
      when 9487 => pixel <= "000000";
      when 9488 => pixel <= "000000";
      when 9489 => pixel <= "000000";
      when 9490 => pixel <= "000000";
      when 9491 => pixel <= "000000";
      when 9492 => pixel <= "001101";
      when 9493 => pixel <= "001101";
      when 9494 => pixel <= "000000";
      when 9495 => pixel <= "000000";
      when 9496 => pixel <= "000000";
      when 9497 => pixel <= "001101";
      when 9498 => pixel <= "001101";
      when 9499 => pixel <= "000000";
      when 9500 => pixel <= "000000";
      when 9501 => pixel <= "000000";
      when 9502 => pixel <= "000000";
      when 9503 => pixel <= "001101";
      when 9504 => pixel <= "001101";
      when 9505 => pixel <= "001101";
      when 9506 => pixel <= "001101";
      when 9507 => pixel <= "000000";
      when 9508 => pixel <= "000000";
      when 9509 => pixel <= "000000";
      when 9510 => pixel <= "000000";
      when 9511 => pixel <= "000000";
      when 9512 => pixel <= "000000";
      when 9513 => pixel <= "000000";
      when 9514 => pixel <= "000000";
      when 9515 => pixel <= "000000";
      when 9516 => pixel <= "000000";
      when 9517 => pixel <= "000000";
      when 9518 => pixel <= "000000";
      when 9519 => pixel <= "001101";
      when 9520 => pixel <= "001101";
      when 9521 => pixel <= "001101";
      when 9522 => pixel <= "000000";
      when 9523 => pixel <= "000000";
      when 9524 => pixel <= "000000";
      when 9525 => pixel <= "001101";
      when 9526 => pixel <= "001101";
      when 9527 => pixel <= "000000";
      when 9528 => pixel <= "000000";
      when 9529 => pixel <= "001101";
      when 9530 => pixel <= "001101";
      when 9531 => pixel <= "000000";
      when 9532 => pixel <= "000000";
      when 9533 => pixel <= "000000";
      when 9534 => pixel <= "000000";
      when 9535 => pixel <= "000000";
      when 9536 => pixel <= "000000";
      when 9537 => pixel <= "000000";
      when 9538 => pixel <= "001101";
      when 9539 => pixel <= "001101";
      when 9540 => pixel <= "000000";
      when 9541 => pixel <= "000000";
      when 9542 => pixel <= "000000";
      when 9543 => pixel <= "001101";
      when 9544 => pixel <= "001101";
      when 9545 => pixel <= "000000";
      when 9546 => pixel <= "000000";
      when 9547 => pixel <= "000000";
      when 9548 => pixel <= "000000";
      when 9549 => pixel <= "000000";
      when 9550 => pixel <= "001101";
      when 9551 => pixel <= "001101";
      when 9552 => pixel <= "000000";
      when 9553 => pixel <= "000000";
      when 9554 => pixel <= "000000";
      when 9555 => pixel <= "000000";
      when 9556 => pixel <= "001101";
      when 9557 => pixel <= "001101";
      when 9558 => pixel <= "000000";
      when 9559 => pixel <= "001101";
      when 9560 => pixel <= "001101";
      when 9561 => pixel <= "001101";
      when 9562 => pixel <= "001101";
      when 9563 => pixel <= "000000";
      when 9564 => pixel <= "000000";
      when 9565 => pixel <= "000000";
      when 9566 => pixel <= "000000";
      when 9567 => pixel <= "000000";
      when 9568 => pixel <= "000000";
      when 9569 => pixel <= "000000";
      when 9570 => pixel <= "000000";
      when 9571 => pixel <= "000000";
      when 9572 => pixel <= "000000";
      when 9573 => pixel <= "000000";
      when 9574 => pixel <= "000000";
      when 9575 => pixel <= "000000";
      when 9576 => pixel <= "000000";
      when 9577 => pixel <= "000000";
      when 9578 => pixel <= "000000";
      when 9579 => pixel <= "000000";
      when 9580 => pixel <= "000000";
      when 9581 => pixel <= "000000";
      when 9582 => pixel <= "000000";
      when 9583 => pixel <= "000000";
      when 9584 => pixel <= "000000";
      when 9585 => pixel <= "000000";
      when 9586 => pixel <= "000000";
      when 9587 => pixel <= "000000";
      when 9588 => pixel <= "000000";
      when 9589 => pixel <= "000000";
      when 9590 => pixel <= "000000";
      when 9591 => pixel <= "000000";
      when 9592 => pixel <= "000000";
      when 9593 => pixel <= "000000";
      when 9594 => pixel <= "000000";
      when 9595 => pixel <= "000000";
      when 9596 => pixel <= "000000";
      when 9597 => pixel <= "000000";
      when 9598 => pixel <= "000000";
      when 9599 => pixel <= "000000";
      when 9600 => pixel <= "000000";
      when 9601 => pixel <= "000000";
      when 9602 => pixel <= "000000";
      when 9603 => pixel <= "000000";
      when 9604 => pixel <= "000000";
      when 9605 => pixel <= "000000";
      when 9606 => pixel <= "000000";
      when 9607 => pixel <= "000000";
      when 9608 => pixel <= "000000";
      when 9609 => pixel <= "000000";
      when 9610 => pixel <= "000000";
      when 9611 => pixel <= "000000";
      when 9612 => pixel <= "000000";
      when 9613 => pixel <= "000000";
      when 9614 => pixel <= "000000";
      when 9615 => pixel <= "000000";
      when 9616 => pixel <= "000000";
      when 9617 => pixel <= "000000";
      when 9618 => pixel <= "000000";
      when 9619 => pixel <= "000000";
      when 9620 => pixel <= "000000";
      when 9621 => pixel <= "000000";
      when 9622 => pixel <= "000000";
      when 9623 => pixel <= "000000";
      when 9624 => pixel <= "000000";
      when 9625 => pixel <= "000000";
      when 9626 => pixel <= "000000";
      when 9627 => pixel <= "000000";
      when 9628 => pixel <= "000000";
      when 9629 => pixel <= "000000";
      when 9630 => pixel <= "000000";
      when 9631 => pixel <= "000000";
      when 9632 => pixel <= "000000";
      when 9633 => pixel <= "000000";
      when 9634 => pixel <= "000000";
      when 9635 => pixel <= "001101";
      when 9636 => pixel <= "001101";
      when 9637 => pixel <= "000000";
      when 9638 => pixel <= "000000";
      when 9639 => pixel <= "000000";
      when 9640 => pixel <= "000000";
      when 9641 => pixel <= "000000";
      when 9642 => pixel <= "000000";
      when 9643 => pixel <= "000000";
      when 9644 => pixel <= "001101";
      when 9645 => pixel <= "001101";
      when 9646 => pixel <= "000000";
      when 9647 => pixel <= "000000";
      when 9648 => pixel <= "000000";
      when 9649 => pixel <= "000000";
      when 9650 => pixel <= "000000";
      when 9651 => pixel <= "000000";
      when 9652 => pixel <= "001101";
      when 9653 => pixel <= "001101";
      when 9654 => pixel <= "001101";
      when 9655 => pixel <= "001101";
      when 9656 => pixel <= "001101";
      when 9657 => pixel <= "001101";
      when 9658 => pixel <= "001101";
      when 9659 => pixel <= "000000";
      when 9660 => pixel <= "000000";
      when 9661 => pixel <= "000000";
      when 9662 => pixel <= "000000";
      when 9663 => pixel <= "000000";
      when 9664 => pixel <= "001101";
      when 9665 => pixel <= "001101";
      when 9666 => pixel <= "000000";
      when 9667 => pixel <= "000000";
      when 9668 => pixel <= "000000";
      when 9669 => pixel <= "000000";
      when 9670 => pixel <= "000000";
      when 9671 => pixel <= "000000";
      when 9672 => pixel <= "000000";
      when 9673 => pixel <= "000000";
      when 9674 => pixel <= "000000";
      when 9675 => pixel <= "000000";
      when 9676 => pixel <= "000000";
      when 9677 => pixel <= "000000";
      when 9678 => pixel <= "000000";
      when 9679 => pixel <= "001101";
      when 9680 => pixel <= "001101";
      when 9681 => pixel <= "001101";
      when 9682 => pixel <= "001101";
      when 9683 => pixel <= "001101";
      when 9684 => pixel <= "001101";
      when 9685 => pixel <= "001101";
      when 9686 => pixel <= "001101";
      when 9687 => pixel <= "000000";
      when 9688 => pixel <= "000000";
      when 9689 => pixel <= "001101";
      when 9690 => pixel <= "001101";
      when 9691 => pixel <= "000000";
      when 9692 => pixel <= "001101";
      when 9693 => pixel <= "001101";
      when 9694 => pixel <= "001101";
      when 9695 => pixel <= "001101";
      when 9696 => pixel <= "000000";
      when 9697 => pixel <= "000000";
      when 9698 => pixel <= "001101";
      when 9699 => pixel <= "001101";
      when 9700 => pixel <= "001101";
      when 9701 => pixel <= "001101";
      when 9702 => pixel <= "001101";
      when 9703 => pixel <= "001101";
      when 9704 => pixel <= "001101";
      when 9705 => pixel <= "000000";
      when 9706 => pixel <= "000000";
      when 9707 => pixel <= "000000";
      when 9708 => pixel <= "000000";
      when 9709 => pixel <= "000000";
      when 9710 => pixel <= "001101";
      when 9711 => pixel <= "001101";
      when 9712 => pixel <= "000000";
      when 9713 => pixel <= "000000";
      when 9714 => pixel <= "000000";
      when 9715 => pixel <= "000000";
      when 9716 => pixel <= "001101";
      when 9717 => pixel <= "001101";
      when 9718 => pixel <= "000000";
      when 9719 => pixel <= "000000";
      when 9720 => pixel <= "001101";
      when 9721 => pixel <= "001101";
      when 9722 => pixel <= "001101";
      when 9723 => pixel <= "000000";
      when 9724 => pixel <= "000000";
      when 9725 => pixel <= "000000";
      when 9726 => pixel <= "000000";
      when 9727 => pixel <= "000000";
      when 9728 => pixel <= "000000";
      when 9729 => pixel <= "000000";
      when 9730 => pixel <= "000000";
      when 9731 => pixel <= "000000";
      when 9732 => pixel <= "000000";
      when 9733 => pixel <= "000000";
      when 9734 => pixel <= "000000";
      when 9735 => pixel <= "000000";
      when 9736 => pixel <= "000000";
      when 9737 => pixel <= "000000";
      when 9738 => pixel <= "000000";
      when 9739 => pixel <= "000000";
      when 9740 => pixel <= "000000";
      when 9741 => pixel <= "000000";
      when 9742 => pixel <= "000000";
      when 9743 => pixel <= "000000";
      when 9744 => pixel <= "000000";
      when 9745 => pixel <= "000000";
      when 9746 => pixel <= "000000";
      when 9747 => pixel <= "000000";
      when 9748 => pixel <= "000000";
      when 9749 => pixel <= "000000";
      when 9750 => pixel <= "000000";
      when 9751 => pixel <= "000000";
      when 9752 => pixel <= "000000";
      when 9753 => pixel <= "000000";
      when 9754 => pixel <= "000000";
      when 9755 => pixel <= "000000";
      when 9756 => pixel <= "000000";
      when 9757 => pixel <= "000000";
      when 9758 => pixel <= "000000";
      when 9759 => pixel <= "000000";
      when 9760 => pixel <= "000000";
      when 9761 => pixel <= "000000";
      when 9762 => pixel <= "000000";
      when 9763 => pixel <= "000000";
      when 9764 => pixel <= "000000";
      when 9765 => pixel <= "000000";
      when 9766 => pixel <= "000000";
      when 9767 => pixel <= "000000";
      when 9768 => pixel <= "000000";
      when 9769 => pixel <= "000000";
      when 9770 => pixel <= "000000";
      when 9771 => pixel <= "000000";
      when 9772 => pixel <= "000000";
      when 9773 => pixel <= "000000";
      when 9774 => pixel <= "000000";
      when 9775 => pixel <= "000000";
      when 9776 => pixel <= "000000";
      when 9777 => pixel <= "000000";
      when 9778 => pixel <= "000000";
      when 9779 => pixel <= "000000";
      when 9780 => pixel <= "000000";
      when 9781 => pixel <= "000000";
      when 9782 => pixel <= "000000";
      when 9783 => pixel <= "000000";
      when 9784 => pixel <= "000000";
      when 9785 => pixel <= "000000";
      when 9786 => pixel <= "000000";
      when 9787 => pixel <= "000000";
      when 9788 => pixel <= "000000";
      when 9789 => pixel <= "000000";
      when 9790 => pixel <= "000000";
      when 9791 => pixel <= "000000";
      when 9792 => pixel <= "000000";
      when 9793 => pixel <= "000000";
      when 9794 => pixel <= "000000";
      when 9795 => pixel <= "001101";
      when 9796 => pixel <= "001101";
      when 9797 => pixel <= "000000";
      when 9798 => pixel <= "000000";
      when 9799 => pixel <= "000000";
      when 9800 => pixel <= "000000";
      when 9801 => pixel <= "000000";
      when 9802 => pixel <= "000000";
      when 9803 => pixel <= "000000";
      when 9804 => pixel <= "001101";
      when 9805 => pixel <= "001101";
      when 9806 => pixel <= "000000";
      when 9807 => pixel <= "000000";
      when 9808 => pixel <= "000000";
      when 9809 => pixel <= "000000";
      when 9810 => pixel <= "000000";
      when 9811 => pixel <= "000000";
      when 9812 => pixel <= "001101";
      when 9813 => pixel <= "001101";
      when 9814 => pixel <= "000000";
      when 9815 => pixel <= "000000";
      when 9816 => pixel <= "000000";
      when 9817 => pixel <= "001101";
      when 9818 => pixel <= "001101";
      when 9819 => pixel <= "000000";
      when 9820 => pixel <= "000000";
      when 9821 => pixel <= "000000";
      when 9822 => pixel <= "000000";
      when 9823 => pixel <= "000000";
      when 9824 => pixel <= "001101";
      when 9825 => pixel <= "001101";
      when 9826 => pixel <= "000000";
      when 9827 => pixel <= "000000";
      when 9828 => pixel <= "000000";
      when 9829 => pixel <= "000000";
      when 9830 => pixel <= "000000";
      when 9831 => pixel <= "000000";
      when 9832 => pixel <= "000000";
      when 9833 => pixel <= "000000";
      when 9834 => pixel <= "000000";
      when 9835 => pixel <= "000000";
      when 9836 => pixel <= "000000";
      when 9837 => pixel <= "000000";
      when 9838 => pixel <= "000000";
      when 9839 => pixel <= "001101";
      when 9840 => pixel <= "001101";
      when 9841 => pixel <= "001101";
      when 9842 => pixel <= "000000";
      when 9843 => pixel <= "000000";
      when 9844 => pixel <= "000000";
      when 9845 => pixel <= "001101";
      when 9846 => pixel <= "001101";
      when 9847 => pixel <= "000000";
      when 9848 => pixel <= "000000";
      when 9849 => pixel <= "001101";
      when 9850 => pixel <= "001101";
      when 9851 => pixel <= "000000";
      when 9852 => pixel <= "000000";
      when 9853 => pixel <= "000000";
      when 9854 => pixel <= "001101";
      when 9855 => pixel <= "001101";
      when 9856 => pixel <= "000000";
      when 9857 => pixel <= "000000";
      when 9858 => pixel <= "001101";
      when 9859 => pixel <= "001101";
      when 9860 => pixel <= "000000";
      when 9861 => pixel <= "000000";
      when 9862 => pixel <= "000000";
      when 9863 => pixel <= "001101";
      when 9864 => pixel <= "001101";
      when 9865 => pixel <= "000000";
      when 9866 => pixel <= "000000";
      when 9867 => pixel <= "000000";
      when 9868 => pixel <= "000000";
      when 9869 => pixel <= "000000";
      when 9870 => pixel <= "001101";
      when 9871 => pixel <= "001101";
      when 9872 => pixel <= "000000";
      when 9873 => pixel <= "000000";
      when 9874 => pixel <= "000000";
      when 9875 => pixel <= "000000";
      when 9876 => pixel <= "001101";
      when 9877 => pixel <= "001101";
      when 9878 => pixel <= "000000";
      when 9879 => pixel <= "000000";
      when 9880 => pixel <= "000000";
      when 9881 => pixel <= "001101";
      when 9882 => pixel <= "001101";
      when 9883 => pixel <= "000000";
      when 9884 => pixel <= "000000";
      when 9885 => pixel <= "000000";
      when 9886 => pixel <= "000000";
      when 9887 => pixel <= "000000";
      when 9888 => pixel <= "000000";
      when 9889 => pixel <= "000000";
      when 9890 => pixel <= "000000";
      when 9891 => pixel <= "000000";
      when 9892 => pixel <= "000000";
      when 9893 => pixel <= "000000";
      when 9894 => pixel <= "000000";
      when 9895 => pixel <= "000000";
      when 9896 => pixel <= "000000";
      when 9897 => pixel <= "000000";
      when 9898 => pixel <= "000000";
      when 9899 => pixel <= "000000";
      when 9900 => pixel <= "000000";
      when 9901 => pixel <= "000000";
      when 9902 => pixel <= "000000";
      when 9903 => pixel <= "000000";
      when 9904 => pixel <= "000000";
      when 9905 => pixel <= "000000";
      when 9906 => pixel <= "000000";
      when 9907 => pixel <= "000000";
      when 9908 => pixel <= "000000";
      when 9909 => pixel <= "000000";
      when 9910 => pixel <= "000000";
      when 9911 => pixel <= "000000";
      when 9912 => pixel <= "000000";
      when 9913 => pixel <= "000000";
      when 9914 => pixel <= "000000";
      when 9915 => pixel <= "000000";
      when 9916 => pixel <= "000000";
      when 9917 => pixel <= "000000";
      when 9918 => pixel <= "000000";
      when 9919 => pixel <= "000000";
      when 9920 => pixel <= "000000";
      when 9921 => pixel <= "000000";
      when 9922 => pixel <= "000000";
      when 9923 => pixel <= "000000";
      when 9924 => pixel <= "000000";
      when 9925 => pixel <= "000000";
      when 9926 => pixel <= "000000";
      when 9927 => pixel <= "000000";
      when 9928 => pixel <= "000000";
      when 9929 => pixel <= "000000";
      when 9930 => pixel <= "000000";
      when 9931 => pixel <= "000000";
      when 9932 => pixel <= "000000";
      when 9933 => pixel <= "000000";
      when 9934 => pixel <= "000000";
      when 9935 => pixel <= "000000";
      when 9936 => pixel <= "000000";
      when 9937 => pixel <= "000000";
      when 9938 => pixel <= "000000";
      when 9939 => pixel <= "000000";
      when 9940 => pixel <= "000000";
      when 9941 => pixel <= "000000";
      when 9942 => pixel <= "000000";
      when 9943 => pixel <= "000000";
      when 9944 => pixel <= "000000";
      when 9945 => pixel <= "000000";
      when 9946 => pixel <= "000000";
      when 9947 => pixel <= "000000";
      when 9948 => pixel <= "000000";
      when 9949 => pixel <= "000000";
      when 9950 => pixel <= "000000";
      when 9951 => pixel <= "000000";
      when 9952 => pixel <= "000000";
      when 9953 => pixel <= "000000";
      when 9954 => pixel <= "000000";
      when 9955 => pixel <= "001101";
      when 9956 => pixel <= "001101";
      when 9957 => pixel <= "000000";
      when 9958 => pixel <= "000000";
      when 9959 => pixel <= "000000";
      when 9960 => pixel <= "000000";
      when 9961 => pixel <= "000000";
      when 9962 => pixel <= "000000";
      when 9963 => pixel <= "000000";
      when 9964 => pixel <= "001101";
      when 9965 => pixel <= "001101";
      when 9966 => pixel <= "000000";
      when 9967 => pixel <= "000000";
      when 9968 => pixel <= "000000";
      when 9969 => pixel <= "001101";
      when 9970 => pixel <= "000000";
      when 9971 => pixel <= "000000";
      when 9972 => pixel <= "001101";
      when 9973 => pixel <= "001101";
      when 9974 => pixel <= "000000";
      when 9975 => pixel <= "000000";
      when 9976 => pixel <= "000000";
      when 9977 => pixel <= "001101";
      when 9978 => pixel <= "001101";
      when 9979 => pixel <= "000000";
      when 9980 => pixel <= "000000";
      when 9981 => pixel <= "000000";
      when 9982 => pixel <= "000000";
      when 9983 => pixel <= "000000";
      when 9984 => pixel <= "001101";
      when 9985 => pixel <= "001101";
      when 9986 => pixel <= "000000";
      when 9987 => pixel <= "000000";
      when 9988 => pixel <= "000000";
      when 9989 => pixel <= "000000";
      when 9990 => pixel <= "000000";
      when 9991 => pixel <= "000000";
      when 9992 => pixel <= "000000";
      when 9993 => pixel <= "000000";
      when 9994 => pixel <= "000000";
      when 9995 => pixel <= "000000";
      when 9996 => pixel <= "000000";
      when 9997 => pixel <= "000000";
      when 9998 => pixel <= "000000";
      when 9999 => pixel <= "001101";
      when 10000 => pixel <= "001101";
      when 10001 => pixel <= "001101";
      when 10002 => pixel <= "000000";
      when 10003 => pixel <= "000000";
      when 10004 => pixel <= "000000";
      when 10005 => pixel <= "001101";
      when 10006 => pixel <= "001101";
      when 10007 => pixel <= "000000";
      when 10008 => pixel <= "000000";
      when 10009 => pixel <= "001101";
      when 10010 => pixel <= "001101";
      when 10011 => pixel <= "000000";
      when 10012 => pixel <= "000000";
      when 10013 => pixel <= "000000";
      when 10014 => pixel <= "001101";
      when 10015 => pixel <= "001101";
      when 10016 => pixel <= "000000";
      when 10017 => pixel <= "000000";
      when 10018 => pixel <= "001101";
      when 10019 => pixel <= "001101";
      when 10020 => pixel <= "000000";
      when 10021 => pixel <= "000000";
      when 10022 => pixel <= "000000";
      when 10023 => pixel <= "001101";
      when 10024 => pixel <= "001101";
      when 10025 => pixel <= "000000";
      when 10026 => pixel <= "000000";
      when 10027 => pixel <= "000000";
      when 10028 => pixel <= "000000";
      when 10029 => pixel <= "000000";
      when 10030 => pixel <= "001101";
      when 10031 => pixel <= "001101";
      when 10032 => pixel <= "000000";
      when 10033 => pixel <= "000000";
      when 10034 => pixel <= "000000";
      when 10035 => pixel <= "000000";
      when 10036 => pixel <= "001101";
      when 10037 => pixel <= "001101";
      when 10038 => pixel <= "000000";
      when 10039 => pixel <= "000000";
      when 10040 => pixel <= "000000";
      when 10041 => pixel <= "001101";
      when 10042 => pixel <= "001101";
      when 10043 => pixel <= "000000";
      when 10044 => pixel <= "000000";
      when 10045 => pixel <= "000000";
      when 10046 => pixel <= "000000";
      when 10047 => pixel <= "000000";
      when 10048 => pixel <= "000000";
      when 10049 => pixel <= "000000";
      when 10050 => pixel <= "000000";
      when 10051 => pixel <= "000000";
      when 10052 => pixel <= "000000";
      when 10053 => pixel <= "000000";
      when 10054 => pixel <= "000000";
      when 10055 => pixel <= "000000";
      when 10056 => pixel <= "000000";
      when 10057 => pixel <= "000000";
      when 10058 => pixel <= "000000";
      when 10059 => pixel <= "000000";
      when 10060 => pixel <= "000000";
      when 10061 => pixel <= "000000";
      when 10062 => pixel <= "000000";
      when 10063 => pixel <= "000000";
      when 10064 => pixel <= "000000";
      when 10065 => pixel <= "000000";
      when 10066 => pixel <= "000000";
      when 10067 => pixel <= "000000";
      when 10068 => pixel <= "000000";
      when 10069 => pixel <= "000000";
      when 10070 => pixel <= "000000";
      when 10071 => pixel <= "000000";
      when 10072 => pixel <= "000000";
      when 10073 => pixel <= "000000";
      when 10074 => pixel <= "000000";
      when 10075 => pixel <= "000000";
      when 10076 => pixel <= "000000";
      when 10077 => pixel <= "000000";
      when 10078 => pixel <= "000000";
      when 10079 => pixel <= "000000";
      when 10080 => pixel <= "000000";
      when 10081 => pixel <= "000000";
      when 10082 => pixel <= "000000";
      when 10083 => pixel <= "000000";
      when 10084 => pixel <= "000000";
      when 10085 => pixel <= "000000";
      when 10086 => pixel <= "000000";
      when 10087 => pixel <= "000000";
      when 10088 => pixel <= "000000";
      when 10089 => pixel <= "000000";
      when 10090 => pixel <= "000000";
      when 10091 => pixel <= "000000";
      when 10092 => pixel <= "000000";
      when 10093 => pixel <= "000000";
      when 10094 => pixel <= "000000";
      when 10095 => pixel <= "000000";
      when 10096 => pixel <= "000000";
      when 10097 => pixel <= "000000";
      when 10098 => pixel <= "000000";
      when 10099 => pixel <= "000000";
      when 10100 => pixel <= "000000";
      when 10101 => pixel <= "000000";
      when 10102 => pixel <= "000000";
      when 10103 => pixel <= "000000";
      when 10104 => pixel <= "000000";
      when 10105 => pixel <= "000000";
      when 10106 => pixel <= "000000";
      when 10107 => pixel <= "000000";
      when 10108 => pixel <= "000000";
      when 10109 => pixel <= "000000";
      when 10110 => pixel <= "000000";
      when 10111 => pixel <= "000000";
      when 10112 => pixel <= "000000";
      when 10113 => pixel <= "000000";
      when 10114 => pixel <= "000000";
      when 10115 => pixel <= "001101";
      when 10116 => pixel <= "001101";
      when 10117 => pixel <= "000000";
      when 10118 => pixel <= "000000";
      when 10119 => pixel <= "000000";
      when 10120 => pixel <= "000000";
      when 10121 => pixel <= "000000";
      when 10122 => pixel <= "000000";
      when 10123 => pixel <= "000000";
      when 10124 => pixel <= "001101";
      when 10125 => pixel <= "001101";
      when 10126 => pixel <= "000000";
      when 10127 => pixel <= "000000";
      when 10128 => pixel <= "001101";
      when 10129 => pixel <= "001101";
      when 10130 => pixel <= "000000";
      when 10131 => pixel <= "000000";
      when 10132 => pixel <= "001101";
      when 10133 => pixel <= "001101";
      when 10134 => pixel <= "000000";
      when 10135 => pixel <= "000000";
      when 10136 => pixel <= "000000";
      when 10137 => pixel <= "001101";
      when 10138 => pixel <= "001101";
      when 10139 => pixel <= "000000";
      when 10140 => pixel <= "000000";
      when 10141 => pixel <= "000000";
      when 10142 => pixel <= "000000";
      when 10143 => pixel <= "000000";
      when 10144 => pixel <= "001101";
      when 10145 => pixel <= "001101";
      when 10146 => pixel <= "000000";
      when 10147 => pixel <= "000000";
      when 10148 => pixel <= "000000";
      when 10149 => pixel <= "000000";
      when 10150 => pixel <= "000000";
      when 10151 => pixel <= "000000";
      when 10152 => pixel <= "000000";
      when 10153 => pixel <= "000000";
      when 10154 => pixel <= "000000";
      when 10155 => pixel <= "000000";
      when 10156 => pixel <= "000000";
      when 10157 => pixel <= "000000";
      when 10158 => pixel <= "000000";
      when 10159 => pixel <= "001101";
      when 10160 => pixel <= "001101";
      when 10161 => pixel <= "001101";
      when 10162 => pixel <= "000000";
      when 10163 => pixel <= "000000";
      when 10164 => pixel <= "000000";
      when 10165 => pixel <= "001101";
      when 10166 => pixel <= "001101";
      when 10167 => pixel <= "000000";
      when 10168 => pixel <= "000000";
      when 10169 => pixel <= "000000";
      when 10170 => pixel <= "001101";
      when 10171 => pixel <= "001101";
      when 10172 => pixel <= "000000";
      when 10173 => pixel <= "000000";
      when 10174 => pixel <= "001101";
      when 10175 => pixel <= "001101";
      when 10176 => pixel <= "000000";
      when 10177 => pixel <= "000000";
      when 10178 => pixel <= "001101";
      when 10179 => pixel <= "001101";
      when 10180 => pixel <= "000000";
      when 10181 => pixel <= "000000";
      when 10182 => pixel <= "000000";
      when 10183 => pixel <= "001101";
      when 10184 => pixel <= "001101";
      when 10185 => pixel <= "000000";
      when 10186 => pixel <= "000000";
      when 10187 => pixel <= "000000";
      when 10188 => pixel <= "000000";
      when 10189 => pixel <= "000000";
      when 10190 => pixel <= "001101";
      when 10191 => pixel <= "001101";
      when 10192 => pixel <= "000000";
      when 10193 => pixel <= "000000";
      when 10194 => pixel <= "000000";
      when 10195 => pixel <= "000000";
      when 10196 => pixel <= "001101";
      when 10197 => pixel <= "001101";
      when 10198 => pixel <= "000000";
      when 10199 => pixel <= "000000";
      when 10200 => pixel <= "000000";
      when 10201 => pixel <= "001101";
      when 10202 => pixel <= "001101";
      when 10203 => pixel <= "000000";
      when 10204 => pixel <= "000000";
      when 10205 => pixel <= "000000";
      when 10206 => pixel <= "000000";
      when 10207 => pixel <= "000000";
      when 10208 => pixel <= "000000";
      when 10209 => pixel <= "000000";
      when 10210 => pixel <= "000000";
      when 10211 => pixel <= "000000";
      when 10212 => pixel <= "000000";
      when 10213 => pixel <= "000000";
      when 10214 => pixel <= "000000";
      when 10215 => pixel <= "000000";
      when 10216 => pixel <= "000000";
      when 10217 => pixel <= "000000";
      when 10218 => pixel <= "000000";
      when 10219 => pixel <= "000000";
      when 10220 => pixel <= "000000";
      when 10221 => pixel <= "000000";
      when 10222 => pixel <= "000000";
      when 10223 => pixel <= "000000";
      when 10224 => pixel <= "000000";
      when 10225 => pixel <= "000000";
      when 10226 => pixel <= "000000";
      when 10227 => pixel <= "000000";
      when 10228 => pixel <= "000000";
      when 10229 => pixel <= "000000";
      when 10230 => pixel <= "000000";
      when 10231 => pixel <= "000000";
      when 10232 => pixel <= "000000";
      when 10233 => pixel <= "000000";
      when 10234 => pixel <= "000000";
      when 10235 => pixel <= "000000";
      when 10236 => pixel <= "000000";
      when 10237 => pixel <= "000000";
      when 10238 => pixel <= "000000";
      when 10239 => pixel <= "000000";
      when 10240 => pixel <= "000000";
      when 10241 => pixel <= "000000";
      when 10242 => pixel <= "000000";
      when 10243 => pixel <= "000000";
      when 10244 => pixel <= "000000";
      when 10245 => pixel <= "000000";
      when 10246 => pixel <= "000000";
      when 10247 => pixel <= "000000";
      when 10248 => pixel <= "000000";
      when 10249 => pixel <= "000000";
      when 10250 => pixel <= "000000";
      when 10251 => pixel <= "000000";
      when 10252 => pixel <= "000000";
      when 10253 => pixel <= "000000";
      when 10254 => pixel <= "000000";
      when 10255 => pixel <= "000000";
      when 10256 => pixel <= "000000";
      when 10257 => pixel <= "000000";
      when 10258 => pixel <= "000000";
      when 10259 => pixel <= "000000";
      when 10260 => pixel <= "000000";
      when 10261 => pixel <= "000000";
      when 10262 => pixel <= "000000";
      when 10263 => pixel <= "000000";
      when 10264 => pixel <= "000000";
      when 10265 => pixel <= "000000";
      when 10266 => pixel <= "000000";
      when 10267 => pixel <= "000000";
      when 10268 => pixel <= "000000";
      when 10269 => pixel <= "000000";
      when 10270 => pixel <= "000000";
      when 10271 => pixel <= "000000";
      when 10272 => pixel <= "000000";
      when 10273 => pixel <= "000000";
      when 10274 => pixel <= "001101";
      when 10275 => pixel <= "001101";
      when 10276 => pixel <= "001101";
      when 10277 => pixel <= "001101";
      when 10278 => pixel <= "000000";
      when 10279 => pixel <= "000000";
      when 10280 => pixel <= "000000";
      when 10281 => pixel <= "000000";
      when 10282 => pixel <= "000000";
      when 10283 => pixel <= "001101";
      when 10284 => pixel <= "001101";
      when 10285 => pixel <= "001101";
      when 10286 => pixel <= "001101";
      when 10287 => pixel <= "001101";
      when 10288 => pixel <= "001101";
      when 10289 => pixel <= "001101";
      when 10290 => pixel <= "000000";
      when 10291 => pixel <= "000000";
      when 10292 => pixel <= "001101";
      when 10293 => pixel <= "001101";
      when 10294 => pixel <= "000000";
      when 10295 => pixel <= "000000";
      when 10296 => pixel <= "000000";
      when 10297 => pixel <= "001101";
      when 10298 => pixel <= "001101";
      when 10299 => pixel <= "000000";
      when 10300 => pixel <= "000000";
      when 10301 => pixel <= "000000";
      when 10302 => pixel <= "000000";
      when 10303 => pixel <= "001101";
      when 10304 => pixel <= "001101";
      when 10305 => pixel <= "001101";
      when 10306 => pixel <= "001101";
      when 10307 => pixel <= "000000";
      when 10308 => pixel <= "000000";
      when 10309 => pixel <= "000000";
      when 10310 => pixel <= "000000";
      when 10311 => pixel <= "000000";
      when 10312 => pixel <= "000000";
      when 10313 => pixel <= "000000";
      when 10314 => pixel <= "000000";
      when 10315 => pixel <= "000000";
      when 10316 => pixel <= "000000";
      when 10317 => pixel <= "000000";
      when 10318 => pixel <= "000000";
      when 10319 => pixel <= "001101";
      when 10320 => pixel <= "001101";
      when 10321 => pixel <= "001101";
      when 10322 => pixel <= "000000";
      when 10323 => pixel <= "000000";
      when 10324 => pixel <= "000000";
      when 10325 => pixel <= "001101";
      when 10326 => pixel <= "001101";
      when 10327 => pixel <= "000000";
      when 10328 => pixel <= "000000";
      when 10329 => pixel <= "000000";
      when 10330 => pixel <= "000000";
      when 10331 => pixel <= "001101";
      when 10332 => pixel <= "001101";
      when 10333 => pixel <= "001101";
      when 10334 => pixel <= "000000";
      when 10335 => pixel <= "001101";
      when 10336 => pixel <= "000000";
      when 10337 => pixel <= "000000";
      when 10338 => pixel <= "001101";
      when 10339 => pixel <= "001101";
      when 10340 => pixel <= "000000";
      when 10341 => pixel <= "000000";
      when 10342 => pixel <= "000000";
      when 10343 => pixel <= "001101";
      when 10344 => pixel <= "001101";
      when 10345 => pixel <= "000000";
      when 10346 => pixel <= "000000";
      when 10347 => pixel <= "000000";
      when 10348 => pixel <= "000000";
      when 10349 => pixel <= "001101";
      when 10350 => pixel <= "001101";
      when 10351 => pixel <= "001101";
      when 10352 => pixel <= "001101";
      when 10353 => pixel <= "000000";
      when 10354 => pixel <= "000000";
      when 10355 => pixel <= "000000";
      when 10356 => pixel <= "001101";
      when 10357 => pixel <= "001101";
      when 10358 => pixel <= "000000";
      when 10359 => pixel <= "000000";
      when 10360 => pixel <= "000000";
      when 10361 => pixel <= "001101";
      when 10362 => pixel <= "001101";
      when 10363 => pixel <= "000000";
      when 10364 => pixel <= "000000";
      when 10365 => pixel <= "000000";
      when 10366 => pixel <= "000000";
      when 10367 => pixel <= "000000";
      when 10368 => pixel <= "000000";
      when 10369 => pixel <= "000000";
      when 10370 => pixel <= "000000";
      when 10371 => pixel <= "000000";
      when 10372 => pixel <= "000000";
      when 10373 => pixel <= "000000";
      when 10374 => pixel <= "000000";
      when 10375 => pixel <= "000000";
      when 10376 => pixel <= "000000";
      when 10377 => pixel <= "000000";
      when 10378 => pixel <= "000000";
      when 10379 => pixel <= "000000";
      when 10380 => pixel <= "000000";
      when 10381 => pixel <= "000000";
      when 10382 => pixel <= "000000";
      when 10383 => pixel <= "000000";
      when 10384 => pixel <= "000000";
      when 10385 => pixel <= "000000";
      when 10386 => pixel <= "000000";
      when 10387 => pixel <= "000000";
      when 10388 => pixel <= "000000";
      when 10389 => pixel <= "000000";
      when 10390 => pixel <= "000000";
      when 10391 => pixel <= "000000";
      when 10392 => pixel <= "000000";
      when 10393 => pixel <= "000000";
      when 10394 => pixel <= "000000";
      when 10395 => pixel <= "000000";
      when 10396 => pixel <= "000000";
      when 10397 => pixel <= "000000";
      when 10398 => pixel <= "000000";
      when 10399 => pixel <= "000000";
      when 10400 => pixel <= "000000";
      when 10401 => pixel <= "000000";
      when 10402 => pixel <= "000000";
      when 10403 => pixel <= "000000";
      when 10404 => pixel <= "000000";
      when 10405 => pixel <= "000000";
      when 10406 => pixel <= "000000";
      when 10407 => pixel <= "000000";
      when 10408 => pixel <= "000000";
      when 10409 => pixel <= "000000";
      when 10410 => pixel <= "000000";
      when 10411 => pixel <= "000000";
      when 10412 => pixel <= "000000";
      when 10413 => pixel <= "000000";
      when 10414 => pixel <= "000000";
      when 10415 => pixel <= "000000";
      when 10416 => pixel <= "000000";
      when 10417 => pixel <= "000000";
      when 10418 => pixel <= "000000";
      when 10419 => pixel <= "000000";
      when 10420 => pixel <= "000000";
      when 10421 => pixel <= "000000";
      when 10422 => pixel <= "000000";
      when 10423 => pixel <= "000000";
      when 10424 => pixel <= "000000";
      when 10425 => pixel <= "000000";
      when 10426 => pixel <= "000000";
      when 10427 => pixel <= "000000";
      when 10428 => pixel <= "000000";
      when 10429 => pixel <= "000000";
      when 10430 => pixel <= "000000";
      when 10431 => pixel <= "000000";
      when 10432 => pixel <= "000000";
      when 10433 => pixel <= "000000";
      when 10434 => pixel <= "000000";
      when 10435 => pixel <= "000000";
      when 10436 => pixel <= "000000";
      when 10437 => pixel <= "000000";
      when 10438 => pixel <= "000000";
      when 10439 => pixel <= "000000";
      when 10440 => pixel <= "000000";
      when 10441 => pixel <= "000000";
      when 10442 => pixel <= "000000";
      when 10443 => pixel <= "000000";
      when 10444 => pixel <= "000000";
      when 10445 => pixel <= "000000";
      when 10446 => pixel <= "000000";
      when 10447 => pixel <= "000000";
      when 10448 => pixel <= "000000";
      when 10449 => pixel <= "000000";
      when 10450 => pixel <= "000000";
      when 10451 => pixel <= "000000";
      when 10452 => pixel <= "000000";
      when 10453 => pixel <= "000000";
      when 10454 => pixel <= "000000";
      when 10455 => pixel <= "000000";
      when 10456 => pixel <= "000000";
      when 10457 => pixel <= "000000";
      when 10458 => pixel <= "000000";
      when 10459 => pixel <= "000000";
      when 10460 => pixel <= "000000";
      when 10461 => pixel <= "000000";
      when 10462 => pixel <= "000000";
      when 10463 => pixel <= "000000";
      when 10464 => pixel <= "000000";
      when 10465 => pixel <= "000000";
      when 10466 => pixel <= "000000";
      when 10467 => pixel <= "000000";
      when 10468 => pixel <= "000000";
      when 10469 => pixel <= "000000";
      when 10470 => pixel <= "000000";
      when 10471 => pixel <= "000000";
      when 10472 => pixel <= "000000";
      when 10473 => pixel <= "000000";
      when 10474 => pixel <= "000000";
      when 10475 => pixel <= "000000";
      when 10476 => pixel <= "000000";
      when 10477 => pixel <= "000000";
      when 10478 => pixel <= "000000";
      when 10479 => pixel <= "000000";
      when 10480 => pixel <= "000000";
      when 10481 => pixel <= "000000";
      when 10482 => pixel <= "000000";
      when 10483 => pixel <= "000000";
      when 10484 => pixel <= "000000";
      when 10485 => pixel <= "000000";
      when 10486 => pixel <= "000000";
      when 10487 => pixel <= "000000";
      when 10488 => pixel <= "000000";
      when 10489 => pixel <= "000000";
      when 10490 => pixel <= "000000";
      when 10491 => pixel <= "000000";
      when 10492 => pixel <= "000000";
      when 10493 => pixel <= "000000";
      when 10494 => pixel <= "000000";
      when 10495 => pixel <= "000000";
      when 10496 => pixel <= "000000";
      when 10497 => pixel <= "000000";
      when 10498 => pixel <= "000000";
      when 10499 => pixel <= "000000";
      when 10500 => pixel <= "000000";
      when 10501 => pixel <= "000000";
      when 10502 => pixel <= "000000";
      when 10503 => pixel <= "000000";
      when 10504 => pixel <= "000000";
      when 10505 => pixel <= "000000";
      when 10506 => pixel <= "000000";
      when 10507 => pixel <= "000000";
      when 10508 => pixel <= "000000";
      when 10509 => pixel <= "000000";
      when 10510 => pixel <= "000000";
      when 10511 => pixel <= "000000";
      when 10512 => pixel <= "000000";
      when 10513 => pixel <= "000000";
      when 10514 => pixel <= "000000";
      when 10515 => pixel <= "000000";
      when 10516 => pixel <= "000000";
      when 10517 => pixel <= "000000";
      when 10518 => pixel <= "000000";
      when 10519 => pixel <= "000000";
      when 10520 => pixel <= "000000";
      when 10521 => pixel <= "000000";
      when 10522 => pixel <= "000000";
      when 10523 => pixel <= "000000";
      when 10524 => pixel <= "000000";
      when 10525 => pixel <= "000000";
      when 10526 => pixel <= "000000";
      when 10527 => pixel <= "000000";
      when 10528 => pixel <= "000000";
      when 10529 => pixel <= "000000";
      when 10530 => pixel <= "000000";
      when 10531 => pixel <= "000000";
      when 10532 => pixel <= "000000";
      when 10533 => pixel <= "000000";
      when 10534 => pixel <= "000000";
      when 10535 => pixel <= "000000";
      when 10536 => pixel <= "000000";
      when 10537 => pixel <= "000000";
      when 10538 => pixel <= "000000";
      when 10539 => pixel <= "000000";
      when 10540 => pixel <= "000000";
      when 10541 => pixel <= "000000";
      when 10542 => pixel <= "000000";
      when 10543 => pixel <= "000000";
      when 10544 => pixel <= "000000";
      when 10545 => pixel <= "000000";
      when 10546 => pixel <= "000000";
      when 10547 => pixel <= "000000";
      when 10548 => pixel <= "000000";
      when 10549 => pixel <= "000000";
      when 10550 => pixel <= "000000";
      when 10551 => pixel <= "000000";
      when 10552 => pixel <= "000000";
      when 10553 => pixel <= "000000";
      when 10554 => pixel <= "000000";
      when 10555 => pixel <= "000000";
      when 10556 => pixel <= "000000";
      when 10557 => pixel <= "000000";
      when 10558 => pixel <= "000000";
      when 10559 => pixel <= "000000";
      when 10560 => pixel <= "000000";
      when 10561 => pixel <= "000000";
      when 10562 => pixel <= "000000";
      when 10563 => pixel <= "000000";
      when 10564 => pixel <= "000000";
      when 10565 => pixel <= "000000";
      when 10566 => pixel <= "000000";
      when 10567 => pixel <= "000000";
      when 10568 => pixel <= "000000";
      when 10569 => pixel <= "000000";
      when 10570 => pixel <= "000000";
      when 10571 => pixel <= "000000";
      when 10572 => pixel <= "000000";
      when 10573 => pixel <= "000000";
      when 10574 => pixel <= "000000";
      when 10575 => pixel <= "000000";
      when 10576 => pixel <= "000000";
      when 10577 => pixel <= "000000";
      when 10578 => pixel <= "000000";
      when 10579 => pixel <= "000000";
      when 10580 => pixel <= "000000";
      when 10581 => pixel <= "000000";
      when 10582 => pixel <= "000000";
      when 10583 => pixel <= "000000";
      when 10584 => pixel <= "000000";
      when 10585 => pixel <= "000000";
      when 10586 => pixel <= "000000";
      when 10587 => pixel <= "000000";
      when 10588 => pixel <= "000000";
      when 10589 => pixel <= "000000";
      when 10590 => pixel <= "000000";
      when 10591 => pixel <= "000000";
      when 10592 => pixel <= "000000";
      when 10593 => pixel <= "000000";
      when 10594 => pixel <= "000000";
      when 10595 => pixel <= "000000";
      when 10596 => pixel <= "000000";
      when 10597 => pixel <= "000000";
      when 10598 => pixel <= "000000";
      when 10599 => pixel <= "000000";
      when 10600 => pixel <= "000000";
      when 10601 => pixel <= "000000";
      when 10602 => pixel <= "000000";
      when 10603 => pixel <= "000000";
      when 10604 => pixel <= "000000";
      when 10605 => pixel <= "000000";
      when 10606 => pixel <= "000000";
      when 10607 => pixel <= "000000";
      when 10608 => pixel <= "000000";
      when 10609 => pixel <= "000000";
      when 10610 => pixel <= "000000";
      when 10611 => pixel <= "000000";
      when 10612 => pixel <= "000000";
      when 10613 => pixel <= "000000";
      when 10614 => pixel <= "000000";
      when 10615 => pixel <= "000000";
      when 10616 => pixel <= "000000";
      when 10617 => pixel <= "000000";
      when 10618 => pixel <= "000000";
      when 10619 => pixel <= "000000";
      when 10620 => pixel <= "000000";
      when 10621 => pixel <= "000000";
      when 10622 => pixel <= "000000";
      when 10623 => pixel <= "000000";
      when 10624 => pixel <= "000000";
      when 10625 => pixel <= "000000";
      when 10626 => pixel <= "000000";
      when 10627 => pixel <= "000000";
      when 10628 => pixel <= "000000";
      when 10629 => pixel <= "000000";
      when 10630 => pixel <= "000000";
      when 10631 => pixel <= "000000";
      when 10632 => pixel <= "000000";
      when 10633 => pixel <= "000000";
      when 10634 => pixel <= "000000";
      when 10635 => pixel <= "000000";
      when 10636 => pixel <= "000000";
      when 10637 => pixel <= "000000";
      when 10638 => pixel <= "000000";
      when 10639 => pixel <= "000000";
      when 10640 => pixel <= "000000";
      when 10641 => pixel <= "000000";
      when 10642 => pixel <= "000000";
      when 10643 => pixel <= "000000";
      when 10644 => pixel <= "000000";
      when 10645 => pixel <= "000000";
      when 10646 => pixel <= "000000";
      when 10647 => pixel <= "000000";
      when 10648 => pixel <= "000000";
      when 10649 => pixel <= "000000";
      when 10650 => pixel <= "000000";
      when 10651 => pixel <= "000000";
      when 10652 => pixel <= "000000";
      when 10653 => pixel <= "000000";
      when 10654 => pixel <= "000000";
      when 10655 => pixel <= "000000";
      when 10656 => pixel <= "000000";
      when 10657 => pixel <= "000000";
      when 10658 => pixel <= "000000";
      when 10659 => pixel <= "000000";
      when 10660 => pixel <= "000000";
      when 10661 => pixel <= "000000";
      when 10662 => pixel <= "000000";
      when 10663 => pixel <= "000000";
      when 10664 => pixel <= "000000";
      when 10665 => pixel <= "000000";
      when 10666 => pixel <= "000000";
      when 10667 => pixel <= "000000";
      when 10668 => pixel <= "000000";
      when 10669 => pixel <= "000000";
      when 10670 => pixel <= "000000";
      when 10671 => pixel <= "000000";
      when 10672 => pixel <= "000000";
      when 10673 => pixel <= "000000";
      when 10674 => pixel <= "000000";
      when 10675 => pixel <= "000000";
      when 10676 => pixel <= "000000";
      when 10677 => pixel <= "000000";
      when 10678 => pixel <= "000000";
      when 10679 => pixel <= "000000";
      when 10680 => pixel <= "000000";
      when 10681 => pixel <= "000000";
      when 10682 => pixel <= "000000";
      when 10683 => pixel <= "000000";
      when 10684 => pixel <= "000000";
      when 10685 => pixel <= "000000";
      when 10686 => pixel <= "000000";
      when 10687 => pixel <= "000000";
      when 10688 => pixel <= "000000";
      when 10689 => pixel <= "000000";
      when 10690 => pixel <= "000000";
      when 10691 => pixel <= "000000";
      when 10692 => pixel <= "000000";
      when 10693 => pixel <= "000000";
      when 10694 => pixel <= "000000";
      when 10695 => pixel <= "000000";
      when 10696 => pixel <= "000000";
      when 10697 => pixel <= "000000";
      when 10698 => pixel <= "000000";
      when 10699 => pixel <= "000000";
      when 10700 => pixel <= "000000";
      when 10701 => pixel <= "000000";
      when 10702 => pixel <= "000000";
      when 10703 => pixel <= "000000";
      when 10704 => pixel <= "000000";
      when 10705 => pixel <= "000000";
      when 10706 => pixel <= "000000";
      when 10707 => pixel <= "000000";
      when 10708 => pixel <= "000000";
      when 10709 => pixel <= "000000";
      when 10710 => pixel <= "000000";
      when 10711 => pixel <= "000000";
      when 10712 => pixel <= "000000";
      when 10713 => pixel <= "000000";
      when 10714 => pixel <= "000000";
      when 10715 => pixel <= "000000";
      when 10716 => pixel <= "000000";
      when 10717 => pixel <= "000000";
      when 10718 => pixel <= "000000";
      when 10719 => pixel <= "000000";
      when 10720 => pixel <= "000000";
      when 10721 => pixel <= "000000";
      when 10722 => pixel <= "000000";
      when 10723 => pixel <= "000000";
      when 10724 => pixel <= "000000";
      when 10725 => pixel <= "000000";
      when 10726 => pixel <= "000000";
      when 10727 => pixel <= "000000";
      when 10728 => pixel <= "000000";
      when 10729 => pixel <= "000000";
      when 10730 => pixel <= "000000";
      when 10731 => pixel <= "000000";
      when 10732 => pixel <= "000000";
      when 10733 => pixel <= "000000";
      when 10734 => pixel <= "000000";
      when 10735 => pixel <= "000000";
      when 10736 => pixel <= "000000";
      when 10737 => pixel <= "000000";
      when 10738 => pixel <= "000000";
      when 10739 => pixel <= "000000";
      when 10740 => pixel <= "000000";
      when 10741 => pixel <= "000000";
      when 10742 => pixel <= "000000";
      when 10743 => pixel <= "000000";
      when 10744 => pixel <= "000000";
      when 10745 => pixel <= "000000";
      when 10746 => pixel <= "000000";
      when 10747 => pixel <= "000000";
      when 10748 => pixel <= "000000";
      when 10749 => pixel <= "000000";
      when 10750 => pixel <= "000000";
      when 10751 => pixel <= "000000";
      when 10752 => pixel <= "000000";
      when 10753 => pixel <= "000000";
      when 10754 => pixel <= "000000";
      when 10755 => pixel <= "000000";
      when 10756 => pixel <= "000000";
      when 10757 => pixel <= "000000";
      when 10758 => pixel <= "000000";
      when 10759 => pixel <= "000000";
      when 10760 => pixel <= "000000";
      when 10761 => pixel <= "000000";
      when 10762 => pixel <= "000000";
      when 10763 => pixel <= "000000";
      when 10764 => pixel <= "000000";
      when 10765 => pixel <= "000000";
      when 10766 => pixel <= "000000";
      when 10767 => pixel <= "000000";
      when 10768 => pixel <= "000000";
      when 10769 => pixel <= "000000";
      when 10770 => pixel <= "000000";
      when 10771 => pixel <= "000000";
      when 10772 => pixel <= "000000";
      when 10773 => pixel <= "000000";
      when 10774 => pixel <= "000000";
      when 10775 => pixel <= "000000";
      when 10776 => pixel <= "000000";
      when 10777 => pixel <= "000000";
      when 10778 => pixel <= "000000";
      when 10779 => pixel <= "000000";
      when 10780 => pixel <= "000000";
      when 10781 => pixel <= "000000";
      when 10782 => pixel <= "000000";
      when 10783 => pixel <= "000000";
      when 10784 => pixel <= "000000";
      when 10785 => pixel <= "000000";
      when 10786 => pixel <= "000000";
      when 10787 => pixel <= "000000";
      when 10788 => pixel <= "000000";
      when 10789 => pixel <= "000000";
      when 10790 => pixel <= "000000";
      when 10791 => pixel <= "000000";
      when 10792 => pixel <= "000000";
      when 10793 => pixel <= "000000";
      when 10794 => pixel <= "000000";
      when 10795 => pixel <= "000000";
      when 10796 => pixel <= "000000";
      when 10797 => pixel <= "000000";
      when 10798 => pixel <= "000000";
      when 10799 => pixel <= "000000";
      when 10800 => pixel <= "000000";
      when 10801 => pixel <= "000000";
      when 10802 => pixel <= "000000";
      when 10803 => pixel <= "000000";
      when 10804 => pixel <= "000000";
      when 10805 => pixel <= "000000";
      when 10806 => pixel <= "000000";
      when 10807 => pixel <= "000000";
      when 10808 => pixel <= "000000";
      when 10809 => pixel <= "000000";
      when 10810 => pixel <= "000000";
      when 10811 => pixel <= "000000";
      when 10812 => pixel <= "000000";
      when 10813 => pixel <= "000000";
      when 10814 => pixel <= "000000";
      when 10815 => pixel <= "000000";
      when 10816 => pixel <= "000000";
      when 10817 => pixel <= "000000";
      when 10818 => pixel <= "000000";
      when 10819 => pixel <= "000000";
      when 10820 => pixel <= "000000";
      when 10821 => pixel <= "000000";
      when 10822 => pixel <= "000000";
      when 10823 => pixel <= "000000";
      when 10824 => pixel <= "000000";
      when 10825 => pixel <= "000000";
      when 10826 => pixel <= "000000";
      when 10827 => pixel <= "000000";
      when 10828 => pixel <= "000000";
      when 10829 => pixel <= "000000";
      when 10830 => pixel <= "000000";
      when 10831 => pixel <= "000000";
      when 10832 => pixel <= "000000";
      when 10833 => pixel <= "000000";
      when 10834 => pixel <= "000000";
      when 10835 => pixel <= "000000";
      when 10836 => pixel <= "000000";
      when 10837 => pixel <= "000000";
      when 10838 => pixel <= "000000";
      when 10839 => pixel <= "000000";
      when 10840 => pixel <= "000000";
      when 10841 => pixel <= "000000";
      when 10842 => pixel <= "000000";
      when 10843 => pixel <= "000000";
      when 10844 => pixel <= "000000";
      when 10845 => pixel <= "000000";
      when 10846 => pixel <= "000000";
      when 10847 => pixel <= "000000";
      when 10848 => pixel <= "000000";
      when 10849 => pixel <= "000000";
      when 10850 => pixel <= "000000";
      when 10851 => pixel <= "000000";
      when 10852 => pixel <= "000000";
      when 10853 => pixel <= "000000";
      when 10854 => pixel <= "000000";
      when 10855 => pixel <= "000000";
      when 10856 => pixel <= "000000";
      when 10857 => pixel <= "000000";
      when 10858 => pixel <= "000000";
      when 10859 => pixel <= "000000";
      when 10860 => pixel <= "000000";
      when 10861 => pixel <= "000000";
      when 10862 => pixel <= "000000";
      when 10863 => pixel <= "000000";
      when 10864 => pixel <= "000000";
      when 10865 => pixel <= "000000";
      when 10866 => pixel <= "000000";
      when 10867 => pixel <= "000000";
      when 10868 => pixel <= "000000";
      when 10869 => pixel <= "000000";
      when 10870 => pixel <= "000000";
      when 10871 => pixel <= "000000";
      when 10872 => pixel <= "000000";
      when 10873 => pixel <= "000000";
      when 10874 => pixel <= "000000";
      when 10875 => pixel <= "000000";
      when 10876 => pixel <= "000000";
      when 10877 => pixel <= "000000";
      when 10878 => pixel <= "000000";
      when 10879 => pixel <= "000000";
      when 10880 => pixel <= "000000";
      when 10881 => pixel <= "000000";
      when 10882 => pixel <= "000000";
      when 10883 => pixel <= "000000";
      when 10884 => pixel <= "000000";
      when 10885 => pixel <= "000000";
      when 10886 => pixel <= "000000";
      when 10887 => pixel <= "000000";
      when 10888 => pixel <= "000000";
      when 10889 => pixel <= "000000";
      when 10890 => pixel <= "000000";
      when 10891 => pixel <= "000000";
      when 10892 => pixel <= "000000";
      when 10893 => pixel <= "000000";
      when 10894 => pixel <= "000000";
      when 10895 => pixel <= "000000";
      when 10896 => pixel <= "000000";
      when 10897 => pixel <= "000000";
      when 10898 => pixel <= "000000";
      when 10899 => pixel <= "000000";
      when 10900 => pixel <= "000000";
      when 10901 => pixel <= "000000";
      when 10902 => pixel <= "000000";
      when 10903 => pixel <= "000000";
      when 10904 => pixel <= "000000";
      when 10905 => pixel <= "000000";
      when 10906 => pixel <= "000000";
      when 10907 => pixel <= "000000";
      when 10908 => pixel <= "000000";
      when 10909 => pixel <= "000000";
      when 10910 => pixel <= "000000";
      when 10911 => pixel <= "000000";
      when 10912 => pixel <= "000000";
      when 10913 => pixel <= "000000";
      when 10914 => pixel <= "000000";
      when 10915 => pixel <= "000000";
      when 10916 => pixel <= "000000";
      when 10917 => pixel <= "000000";
      when 10918 => pixel <= "000000";
      when 10919 => pixel <= "000000";
      when 10920 => pixel <= "000000";
      when 10921 => pixel <= "000000";
      when 10922 => pixel <= "000000";
      when 10923 => pixel <= "000000";
      when 10924 => pixel <= "000000";
      when 10925 => pixel <= "000000";
      when 10926 => pixel <= "000000";
      when 10927 => pixel <= "000000";
      when 10928 => pixel <= "000000";
      when 10929 => pixel <= "000000";
      when 10930 => pixel <= "000000";
      when 10931 => pixel <= "000000";
      when 10932 => pixel <= "000000";
      when 10933 => pixel <= "000000";
      when 10934 => pixel <= "000000";
      when 10935 => pixel <= "000000";
      when 10936 => pixel <= "000000";
      when 10937 => pixel <= "000000";
      when 10938 => pixel <= "000000";
      when 10939 => pixel <= "000000";
      when 10940 => pixel <= "000000";
      when 10941 => pixel <= "000000";
      when 10942 => pixel <= "000000";
      when 10943 => pixel <= "000000";
      when 10944 => pixel <= "000000";
      when 10945 => pixel <= "000000";
      when 10946 => pixel <= "000000";
      when 10947 => pixel <= "000000";
      when 10948 => pixel <= "000000";
      when 10949 => pixel <= "000000";
      when 10950 => pixel <= "000000";
      when 10951 => pixel <= "000000";
      when 10952 => pixel <= "000000";
      when 10953 => pixel <= "000000";
      when 10954 => pixel <= "000000";
      when 10955 => pixel <= "000000";
      when 10956 => pixel <= "000000";
      when 10957 => pixel <= "000000";
      when 10958 => pixel <= "000000";
      when 10959 => pixel <= "000000";
      when 10960 => pixel <= "000000";
      when 10961 => pixel <= "000000";
      when 10962 => pixel <= "000000";
      when 10963 => pixel <= "000000";
      when 10964 => pixel <= "000000";
      when 10965 => pixel <= "000000";
      when 10966 => pixel <= "000000";
      when 10967 => pixel <= "000000";
      when 10968 => pixel <= "000000";
      when 10969 => pixel <= "000000";
      when 10970 => pixel <= "000000";
      when 10971 => pixel <= "000000";
      when 10972 => pixel <= "000000";
      when 10973 => pixel <= "000000";
      when 10974 => pixel <= "000000";
      when 10975 => pixel <= "000000";
      when 10976 => pixel <= "000000";
      when 10977 => pixel <= "000000";
      when 10978 => pixel <= "000000";
      when 10979 => pixel <= "000000";
      when 10980 => pixel <= "000000";
      when 10981 => pixel <= "000000";
      when 10982 => pixel <= "000000";
      when 10983 => pixel <= "000000";
      when 10984 => pixel <= "000000";
      when 10985 => pixel <= "000000";
      when 10986 => pixel <= "000000";
      when 10987 => pixel <= "000000";
      when 10988 => pixel <= "000000";
      when 10989 => pixel <= "000000";
      when 10990 => pixel <= "000000";
      when 10991 => pixel <= "000000";
      when 10992 => pixel <= "000000";
      when 10993 => pixel <= "000000";
      when 10994 => pixel <= "000000";
      when 10995 => pixel <= "000000";
      when 10996 => pixel <= "000000";
      when 10997 => pixel <= "000000";
      when 10998 => pixel <= "000000";
      when 10999 => pixel <= "000000";
      when 11000 => pixel <= "000000";
      when 11001 => pixel <= "000000";
      when 11002 => pixel <= "000000";
      when 11003 => pixel <= "000000";
      when 11004 => pixel <= "000000";
      when 11005 => pixel <= "000000";
      when 11006 => pixel <= "000000";
      when 11007 => pixel <= "000000";
      when 11008 => pixel <= "000000";
      when 11009 => pixel <= "000000";
      when 11010 => pixel <= "000000";
      when 11011 => pixel <= "000000";
      when 11012 => pixel <= "000000";
      when 11013 => pixel <= "000000";
      when 11014 => pixel <= "000000";
      when 11015 => pixel <= "000000";
      when 11016 => pixel <= "000000";
      when 11017 => pixel <= "000000";
      when 11018 => pixel <= "000000";
      when 11019 => pixel <= "000000";
      when 11020 => pixel <= "000000";
      when 11021 => pixel <= "000000";
      when 11022 => pixel <= "000000";
      when 11023 => pixel <= "000000";
      when 11024 => pixel <= "000000";
      when 11025 => pixel <= "000000";
      when 11026 => pixel <= "000000";
      when 11027 => pixel <= "000000";
      when 11028 => pixel <= "000000";
      when 11029 => pixel <= "000000";
      when 11030 => pixel <= "000000";
      when 11031 => pixel <= "000000";
      when 11032 => pixel <= "000000";
      when 11033 => pixel <= "000000";
      when 11034 => pixel <= "000000";
      when 11035 => pixel <= "000000";
      when 11036 => pixel <= "000000";
      when 11037 => pixel <= "000000";
      when 11038 => pixel <= "000000";
      when 11039 => pixel <= "000000";
      when 11040 => pixel <= "000000";
      when 11041 => pixel <= "000000";
      when 11042 => pixel <= "000000";
      when 11043 => pixel <= "000000";
      when 11044 => pixel <= "000000";
      when 11045 => pixel <= "000000";
      when 11046 => pixel <= "000000";
      when 11047 => pixel <= "000000";
      when 11048 => pixel <= "000000";
      when 11049 => pixel <= "000000";
      when 11050 => pixel <= "000000";
      when 11051 => pixel <= "000000";
      when 11052 => pixel <= "000000";
      when 11053 => pixel <= "000000";
      when 11054 => pixel <= "000000";
      when 11055 => pixel <= "000000";
      when 11056 => pixel <= "000000";
      when 11057 => pixel <= "000000";
      when 11058 => pixel <= "000000";
      when 11059 => pixel <= "000000";
      when 11060 => pixel <= "000000";
      when 11061 => pixel <= "000000";
      when 11062 => pixel <= "000000";
      when 11063 => pixel <= "000000";
      when 11064 => pixel <= "000000";
      when 11065 => pixel <= "000000";
      when 11066 => pixel <= "000000";
      when 11067 => pixel <= "000000";
      when 11068 => pixel <= "000000";
      when 11069 => pixel <= "000000";
      when 11070 => pixel <= "000000";
      when 11071 => pixel <= "000000";
      when 11072 => pixel <= "000000";
      when 11073 => pixel <= "000000";
      when 11074 => pixel <= "000000";
      when 11075 => pixel <= "000000";
      when 11076 => pixel <= "000000";
      when 11077 => pixel <= "000000";
      when 11078 => pixel <= "000000";
      when 11079 => pixel <= "000000";
      when 11080 => pixel <= "000000";
      when 11081 => pixel <= "000000";
      when 11082 => pixel <= "000000";
      when 11083 => pixel <= "000000";
      when 11084 => pixel <= "000000";
      when 11085 => pixel <= "000000";
      when 11086 => pixel <= "000000";
      when 11087 => pixel <= "000000";
      when 11088 => pixel <= "000000";
      when 11089 => pixel <= "000000";
      when 11090 => pixel <= "000000";
      when 11091 => pixel <= "000000";
      when 11092 => pixel <= "000000";
      when 11093 => pixel <= "000000";
      when 11094 => pixel <= "000000";
      when 11095 => pixel <= "000000";
      when 11096 => pixel <= "000000";
      when 11097 => pixel <= "000000";
      when 11098 => pixel <= "000000";
      when 11099 => pixel <= "000000";
      when 11100 => pixel <= "000000";
      when 11101 => pixel <= "000000";
      when 11102 => pixel <= "000000";
      when 11103 => pixel <= "000000";
      when 11104 => pixel <= "000000";
      when 11105 => pixel <= "000000";
      when 11106 => pixel <= "000000";
      when 11107 => pixel <= "000000";
      when 11108 => pixel <= "000000";
      when 11109 => pixel <= "000000";
      when 11110 => pixel <= "000000";
      when 11111 => pixel <= "000000";
      when 11112 => pixel <= "000000";
      when 11113 => pixel <= "000000";
      when 11114 => pixel <= "000000";
      when 11115 => pixel <= "000000";
      when 11116 => pixel <= "000000";
      when 11117 => pixel <= "000000";
      when 11118 => pixel <= "000000";
      when 11119 => pixel <= "000000";
      when 11120 => pixel <= "000000";
      when 11121 => pixel <= "000000";
      when 11122 => pixel <= "000000";
      when 11123 => pixel <= "000000";
      when 11124 => pixel <= "000000";
      when 11125 => pixel <= "000000";
      when 11126 => pixel <= "000000";
      when 11127 => pixel <= "000000";
      when 11128 => pixel <= "000000";
      when 11129 => pixel <= "000000";
      when 11130 => pixel <= "000000";
      when 11131 => pixel <= "000000";
      when 11132 => pixel <= "000000";
      when 11133 => pixel <= "000000";
      when 11134 => pixel <= "000000";
      when 11135 => pixel <= "000000";
      when 11136 => pixel <= "000000";
      when 11137 => pixel <= "000000";
      when 11138 => pixel <= "000000";
      when 11139 => pixel <= "000000";
      when 11140 => pixel <= "000000";
      when 11141 => pixel <= "000000";
      when 11142 => pixel <= "000000";
      when 11143 => pixel <= "000000";
      when 11144 => pixel <= "000000";
      when 11145 => pixel <= "000000";
      when 11146 => pixel <= "000000";
      when 11147 => pixel <= "000000";
      when 11148 => pixel <= "000000";
      when 11149 => pixel <= "000000";
      when 11150 => pixel <= "000000";
      when 11151 => pixel <= "000000";
      when 11152 => pixel <= "000000";
      when 11153 => pixel <= "000000";
      when 11154 => pixel <= "000000";
      when 11155 => pixel <= "000000";
      when 11156 => pixel <= "000000";
      when 11157 => pixel <= "000000";
      when 11158 => pixel <= "000000";
      when 11159 => pixel <= "000000";
      when 11160 => pixel <= "000000";
      when 11161 => pixel <= "000000";
      when 11162 => pixel <= "000000";
      when 11163 => pixel <= "000000";
      when 11164 => pixel <= "000000";
      when 11165 => pixel <= "000000";
      when 11166 => pixel <= "000000";
      when 11167 => pixel <= "000000";
      when 11168 => pixel <= "000000";
      when 11169 => pixel <= "000000";
      when 11170 => pixel <= "000000";
      when 11171 => pixel <= "000000";
      when 11172 => pixel <= "000000";
      when 11173 => pixel <= "000000";
      when 11174 => pixel <= "000000";
      when 11175 => pixel <= "000000";
      when 11176 => pixel <= "000000";
      when 11177 => pixel <= "000000";
      when 11178 => pixel <= "000000";
      when 11179 => pixel <= "000000";
      when 11180 => pixel <= "000000";
      when 11181 => pixel <= "000000";
      when 11182 => pixel <= "000000";
      when 11183 => pixel <= "000000";
      when 11184 => pixel <= "000000";
      when 11185 => pixel <= "000000";
      when 11186 => pixel <= "000000";
      when 11187 => pixel <= "000000";
      when 11188 => pixel <= "000000";
      when 11189 => pixel <= "000000";
      when 11190 => pixel <= "000000";
      when 11191 => pixel <= "000000";
      when 11192 => pixel <= "000000";
      when 11193 => pixel <= "000000";
      when 11194 => pixel <= "000000";
      when 11195 => pixel <= "000000";
      when 11196 => pixel <= "000000";
      when 11197 => pixel <= "000000";
      when 11198 => pixel <= "000000";
      when 11199 => pixel <= "000000";
      when 11200 => pixel <= "000000";
      when 11201 => pixel <= "000000";
      when 11202 => pixel <= "000000";
      when 11203 => pixel <= "000000";
      when 11204 => pixel <= "000000";
      when 11205 => pixel <= "000000";
      when 11206 => pixel <= "000000";
      when 11207 => pixel <= "000000";
      when 11208 => pixel <= "000000";
      when 11209 => pixel <= "000000";
      when 11210 => pixel <= "000000";
      when 11211 => pixel <= "000000";
      when 11212 => pixel <= "000000";
      when 11213 => pixel <= "000000";
      when 11214 => pixel <= "000000";
      when 11215 => pixel <= "000000";
      when 11216 => pixel <= "000000";
      when 11217 => pixel <= "000000";
      when 11218 => pixel <= "000000";
      when 11219 => pixel <= "000000";
      when 11220 => pixel <= "000000";
      when 11221 => pixel <= "000000";
      when 11222 => pixel <= "000000";
      when 11223 => pixel <= "000000";
      when 11224 => pixel <= "000000";
      when 11225 => pixel <= "000000";
      when 11226 => pixel <= "000000";
      when 11227 => pixel <= "000000";
      when 11228 => pixel <= "000000";
      when 11229 => pixel <= "000000";
      when 11230 => pixel <= "000000";
      when 11231 => pixel <= "000000";
      when 11232 => pixel <= "000000";
      when 11233 => pixel <= "000000";
      when 11234 => pixel <= "000000";
      when 11235 => pixel <= "000000";
      when 11236 => pixel <= "000000";
      when 11237 => pixel <= "000000";
      when 11238 => pixel <= "000000";
      when 11239 => pixel <= "000000";
      when 11240 => pixel <= "000000";
      when 11241 => pixel <= "000000";
      when 11242 => pixel <= "000000";
      when 11243 => pixel <= "000000";
      when 11244 => pixel <= "000000";
      when 11245 => pixel <= "000000";
      when 11246 => pixel <= "000000";
      when 11247 => pixel <= "000000";
      when 11248 => pixel <= "000000";
      when 11249 => pixel <= "000000";
      when 11250 => pixel <= "000000";
      when 11251 => pixel <= "000000";
      when 11252 => pixel <= "000000";
      when 11253 => pixel <= "000000";
      when 11254 => pixel <= "000000";
      when 11255 => pixel <= "000000";
      when 11256 => pixel <= "000000";
      when 11257 => pixel <= "000000";
      when 11258 => pixel <= "000000";
      when 11259 => pixel <= "000000";
      when 11260 => pixel <= "000000";
      when 11261 => pixel <= "000000";
      when 11262 => pixel <= "000000";
      when 11263 => pixel <= "000000";
      when 11264 => pixel <= "000000";
      when 11265 => pixel <= "000000";
      when 11266 => pixel <= "000000";
      when 11267 => pixel <= "000000";
      when 11268 => pixel <= "000000";
      when 11269 => pixel <= "000000";
      when 11270 => pixel <= "000000";
      when 11271 => pixel <= "000000";
      when 11272 => pixel <= "000000";
      when 11273 => pixel <= "000000";
      when 11274 => pixel <= "000000";
      when 11275 => pixel <= "000000";
      when 11276 => pixel <= "000000";
      when 11277 => pixel <= "000000";
      when 11278 => pixel <= "000000";
      when 11279 => pixel <= "000000";
      when 11280 => pixel <= "000000";
      when 11281 => pixel <= "000000";
      when 11282 => pixel <= "000000";
      when 11283 => pixel <= "000000";
      when 11284 => pixel <= "000000";
      when 11285 => pixel <= "000000";
      when 11286 => pixel <= "000000";
      when 11287 => pixel <= "000000";
      when 11288 => pixel <= "000000";
      when 11289 => pixel <= "000000";
      when 11290 => pixel <= "000000";
      when 11291 => pixel <= "000000";
      when 11292 => pixel <= "000000";
      when 11293 => pixel <= "000000";
      when 11294 => pixel <= "000000";
      when 11295 => pixel <= "000000";
      when 11296 => pixel <= "000000";
      when 11297 => pixel <= "000000";
      when 11298 => pixel <= "000000";
      when 11299 => pixel <= "000000";
      when 11300 => pixel <= "000000";
      when 11301 => pixel <= "000000";
      when 11302 => pixel <= "000000";
      when 11303 => pixel <= "000000";
      when 11304 => pixel <= "000000";
      when 11305 => pixel <= "000000";
      when 11306 => pixel <= "000000";
      when 11307 => pixel <= "000000";
      when 11308 => pixel <= "000000";
      when 11309 => pixel <= "000000";
      when 11310 => pixel <= "000000";
      when 11311 => pixel <= "000000";
      when 11312 => pixel <= "000000";
      when 11313 => pixel <= "000000";
      when 11314 => pixel <= "000000";
      when 11315 => pixel <= "000000";
      when 11316 => pixel <= "000000";
      when 11317 => pixel <= "000000";
      when 11318 => pixel <= "000000";
      when 11319 => pixel <= "000000";
      when 11320 => pixel <= "000000";
      when 11321 => pixel <= "000000";
      when 11322 => pixel <= "000000";
      when 11323 => pixel <= "000000";
      when 11324 => pixel <= "000000";
      when 11325 => pixel <= "000000";
      when 11326 => pixel <= "000000";
      when 11327 => pixel <= "000000";
      when 11328 => pixel <= "000000";
      when 11329 => pixel <= "000000";
      when 11330 => pixel <= "000000";
      when 11331 => pixel <= "000000";
      when 11332 => pixel <= "000000";
      when 11333 => pixel <= "000000";
      when 11334 => pixel <= "000000";
      when 11335 => pixel <= "000000";
      when 11336 => pixel <= "000000";
      when 11337 => pixel <= "000000";
      when 11338 => pixel <= "000000";
      when 11339 => pixel <= "000000";
      when 11340 => pixel <= "000000";
      when 11341 => pixel <= "000000";
      when 11342 => pixel <= "000000";
      when 11343 => pixel <= "000000";
      when 11344 => pixel <= "000000";
      when 11345 => pixel <= "000000";
      when 11346 => pixel <= "000000";
      when 11347 => pixel <= "000000";
      when 11348 => pixel <= "000000";
      when 11349 => pixel <= "000000";
      when 11350 => pixel <= "000000";
      when 11351 => pixel <= "000000";
      when 11352 => pixel <= "000000";
      when 11353 => pixel <= "000000";
      when 11354 => pixel <= "000000";
      when 11355 => pixel <= "000000";
      when 11356 => pixel <= "000000";
      when 11357 => pixel <= "000000";
      when 11358 => pixel <= "000000";
      when 11359 => pixel <= "000000";
      when 11360 => pixel <= "000000";
      when 11361 => pixel <= "000000";
      when 11362 => pixel <= "000000";
      when 11363 => pixel <= "000000";
      when 11364 => pixel <= "000000";
      when 11365 => pixel <= "000000";
      when 11366 => pixel <= "000000";
      when 11367 => pixel <= "000000";
      when 11368 => pixel <= "000000";
      when 11369 => pixel <= "000000";
      when 11370 => pixel <= "000000";
      when 11371 => pixel <= "000000";
      when 11372 => pixel <= "000000";
      when 11373 => pixel <= "000000";
      when 11374 => pixel <= "000000";
      when 11375 => pixel <= "000000";
      when 11376 => pixel <= "000000";
      when 11377 => pixel <= "000000";
      when 11378 => pixel <= "000000";
      when 11379 => pixel <= "000000";
      when 11380 => pixel <= "000000";
      when 11381 => pixel <= "000000";
      when 11382 => pixel <= "000000";
      when 11383 => pixel <= "000000";
      when 11384 => pixel <= "000000";
      when 11385 => pixel <= "000000";
      when 11386 => pixel <= "000000";
      when 11387 => pixel <= "000000";
      when 11388 => pixel <= "000000";
      when 11389 => pixel <= "000000";
      when 11390 => pixel <= "000000";
      when 11391 => pixel <= "000000";
      when 11392 => pixel <= "000000";
      when 11393 => pixel <= "000000";
      when 11394 => pixel <= "000000";
      when 11395 => pixel <= "000000";
      when 11396 => pixel <= "000000";
      when 11397 => pixel <= "000000";
      when 11398 => pixel <= "000000";
      when 11399 => pixel <= "000000";
      when 11400 => pixel <= "000000";
      when 11401 => pixel <= "000000";
      when 11402 => pixel <= "000000";
      when 11403 => pixel <= "000000";
      when 11404 => pixel <= "000000";
      when 11405 => pixel <= "000000";
      when 11406 => pixel <= "000000";
      when 11407 => pixel <= "000000";
      when 11408 => pixel <= "000000";
      when 11409 => pixel <= "000000";
      when 11410 => pixel <= "000000";
      when 11411 => pixel <= "000000";
      when 11412 => pixel <= "000000";
      when 11413 => pixel <= "000000";
      when 11414 => pixel <= "000000";
      when 11415 => pixel <= "000000";
      when 11416 => pixel <= "000000";
      when 11417 => pixel <= "000000";
      when 11418 => pixel <= "000000";
      when 11419 => pixel <= "000000";
      when 11420 => pixel <= "000000";
      when 11421 => pixel <= "000000";
      when 11422 => pixel <= "000000";
      when 11423 => pixel <= "000000";
      when 11424 => pixel <= "000000";
      when 11425 => pixel <= "000000";
      when 11426 => pixel <= "000000";
      when 11427 => pixel <= "000000";
      when 11428 => pixel <= "000000";
      when 11429 => pixel <= "000000";
      when 11430 => pixel <= "000000";
      when 11431 => pixel <= "000000";
      when 11432 => pixel <= "000000";
      when 11433 => pixel <= "000000";
      when 11434 => pixel <= "000000";
      when 11435 => pixel <= "000000";
      when 11436 => pixel <= "000000";
      when 11437 => pixel <= "000000";
      when 11438 => pixel <= "000000";
      when 11439 => pixel <= "000000";
      when 11440 => pixel <= "000000";
      when 11441 => pixel <= "000000";
      when 11442 => pixel <= "000000";
      when 11443 => pixel <= "000000";
      when 11444 => pixel <= "000000";
      when 11445 => pixel <= "000000";
      when 11446 => pixel <= "000000";
      when 11447 => pixel <= "000000";
      when 11448 => pixel <= "000000";
      when 11449 => pixel <= "000000";
      when 11450 => pixel <= "000000";
      when 11451 => pixel <= "000000";
      when 11452 => pixel <= "000000";
      when 11453 => pixel <= "000000";
      when 11454 => pixel <= "000000";
      when 11455 => pixel <= "000000";
      when 11456 => pixel <= "000000";
      when 11457 => pixel <= "000000";
      when 11458 => pixel <= "000000";
      when 11459 => pixel <= "000000";
      when 11460 => pixel <= "000000";
      when 11461 => pixel <= "000000";
      when 11462 => pixel <= "000000";
      when 11463 => pixel <= "000000";
      when 11464 => pixel <= "000000";
      when 11465 => pixel <= "000000";
      when 11466 => pixel <= "000000";
      when 11467 => pixel <= "000000";
      when 11468 => pixel <= "000000";
      when 11469 => pixel <= "000000";
      when 11470 => pixel <= "000000";
      when 11471 => pixel <= "000000";
      when 11472 => pixel <= "000000";
      when 11473 => pixel <= "000000";
      when 11474 => pixel <= "000000";
      when 11475 => pixel <= "000000";
      when 11476 => pixel <= "000000";
      when 11477 => pixel <= "000000";
      when 11478 => pixel <= "000000";
      when 11479 => pixel <= "000000";
      when 11480 => pixel <= "000000";
      when 11481 => pixel <= "000000";
      when 11482 => pixel <= "000000";
      when 11483 => pixel <= "000000";
      when 11484 => pixel <= "000000";
      when 11485 => pixel <= "000000";
      when 11486 => pixel <= "000000";
      when 11487 => pixel <= "000000";
      when 11488 => pixel <= "000000";
      when 11489 => pixel <= "000000";
      when 11490 => pixel <= "000000";
      when 11491 => pixel <= "000000";
      when 11492 => pixel <= "000000";
      when 11493 => pixel <= "000000";
      when 11494 => pixel <= "000000";
      when 11495 => pixel <= "000000";
      when 11496 => pixel <= "000000";
      when 11497 => pixel <= "000000";
      when 11498 => pixel <= "000000";
      when 11499 => pixel <= "000000";
      when 11500 => pixel <= "000000";
      when 11501 => pixel <= "000000";
      when 11502 => pixel <= "000000";
      when 11503 => pixel <= "000000";
      when 11504 => pixel <= "000000";
      when 11505 => pixel <= "000000";
      when 11506 => pixel <= "000000";
      when 11507 => pixel <= "000000";
      when 11508 => pixel <= "000000";
      when 11509 => pixel <= "000000";
      when 11510 => pixel <= "000000";
      when 11511 => pixel <= "000000";
      when 11512 => pixel <= "000000";
      when 11513 => pixel <= "000000";
      when 11514 => pixel <= "000000";
      when 11515 => pixel <= "000000";
      when 11516 => pixel <= "000000";
      when 11517 => pixel <= "000000";
      when 11518 => pixel <= "000000";
      when 11519 => pixel <= "000000";
      when 11520 => pixel <= "000000";
      when 11521 => pixel <= "000000";
      when 11522 => pixel <= "000000";
      when 11523 => pixel <= "000000";
      when 11524 => pixel <= "000000";
      when 11525 => pixel <= "000000";
      when 11526 => pixel <= "000000";
      when 11527 => pixel <= "000000";
      when 11528 => pixel <= "000000";
      when 11529 => pixel <= "000000";
      when 11530 => pixel <= "000000";
      when 11531 => pixel <= "000000";
      when 11532 => pixel <= "000000";
      when 11533 => pixel <= "000000";
      when 11534 => pixel <= "000000";
      when 11535 => pixel <= "000000";
      when 11536 => pixel <= "000000";
      when 11537 => pixel <= "000000";
      when 11538 => pixel <= "000000";
      when 11539 => pixel <= "000000";
      when 11540 => pixel <= "000000";
      when 11541 => pixel <= "000000";
      when 11542 => pixel <= "000000";
      when 11543 => pixel <= "000000";
      when 11544 => pixel <= "000000";
      when 11545 => pixel <= "000000";
      when 11546 => pixel <= "000000";
      when 11547 => pixel <= "000000";
      when 11548 => pixel <= "000000";
      when 11549 => pixel <= "000000";
      when 11550 => pixel <= "000000";
      when 11551 => pixel <= "000000";
      when 11552 => pixel <= "000000";
      when 11553 => pixel <= "000000";
      when 11554 => pixel <= "000000";
      when 11555 => pixel <= "000000";
      when 11556 => pixel <= "000000";
      when 11557 => pixel <= "000000";
      when 11558 => pixel <= "000000";
      when 11559 => pixel <= "000000";
      when 11560 => pixel <= "000000";
      when 11561 => pixel <= "000000";
      when 11562 => pixel <= "000000";
      when 11563 => pixel <= "000000";
      when 11564 => pixel <= "000000";
      when 11565 => pixel <= "000000";
      when 11566 => pixel <= "000000";
      when 11567 => pixel <= "000000";
      when 11568 => pixel <= "000000";
      when 11569 => pixel <= "000000";
      when 11570 => pixel <= "000000";
      when 11571 => pixel <= "000000";
      when 11572 => pixel <= "000000";
      when 11573 => pixel <= "000000";
      when 11574 => pixel <= "000000";
      when 11575 => pixel <= "000000";
      when 11576 => pixel <= "000000";
      when 11577 => pixel <= "000000";
      when 11578 => pixel <= "000000";
      when 11579 => pixel <= "000000";
      when 11580 => pixel <= "000000";
      when 11581 => pixel <= "000000";
      when 11582 => pixel <= "000000";
      when 11583 => pixel <= "000000";
      when 11584 => pixel <= "000000";
      when 11585 => pixel <= "000000";
      when 11586 => pixel <= "000000";
      when 11587 => pixel <= "000000";
      when 11588 => pixel <= "000000";
      when 11589 => pixel <= "000000";
      when 11590 => pixel <= "000000";
      when 11591 => pixel <= "000000";
      when 11592 => pixel <= "000000";
      when 11593 => pixel <= "000000";
      when 11594 => pixel <= "000000";
      when 11595 => pixel <= "000000";
      when 11596 => pixel <= "000000";
      when 11597 => pixel <= "000000";
      when 11598 => pixel <= "000000";
      when 11599 => pixel <= "000000";
      when 11600 => pixel <= "000000";
      when 11601 => pixel <= "000000";
      when 11602 => pixel <= "000000";
      when 11603 => pixel <= "000000";
      when 11604 => pixel <= "000000";
      when 11605 => pixel <= "000000";
      when 11606 => pixel <= "000000";
      when 11607 => pixel <= "000000";
      when 11608 => pixel <= "000000";
      when 11609 => pixel <= "000000";
      when 11610 => pixel <= "000000";
      when 11611 => pixel <= "000000";
      when 11612 => pixel <= "000000";
      when 11613 => pixel <= "000000";
      when 11614 => pixel <= "000000";
      when 11615 => pixel <= "000000";
      when 11616 => pixel <= "000000";
      when 11617 => pixel <= "000000";
      when 11618 => pixel <= "000000";
      when 11619 => pixel <= "000000";
      when 11620 => pixel <= "000000";
      when 11621 => pixel <= "000000";
      when 11622 => pixel <= "000000";
      when 11623 => pixel <= "000000";
      when 11624 => pixel <= "000000";
      when 11625 => pixel <= "000000";
      when 11626 => pixel <= "000000";
      when 11627 => pixel <= "000000";
      when 11628 => pixel <= "000000";
      when 11629 => pixel <= "000000";
      when 11630 => pixel <= "000000";
      when 11631 => pixel <= "000000";
      when 11632 => pixel <= "000000";
      when 11633 => pixel <= "000000";
      when 11634 => pixel <= "000000";
      when 11635 => pixel <= "000000";
      when 11636 => pixel <= "000000";
      when 11637 => pixel <= "000000";
      when 11638 => pixel <= "000000";
      when 11639 => pixel <= "000000";
      when 11640 => pixel <= "000000";
      when 11641 => pixel <= "000000";
      when 11642 => pixel <= "000000";
      when 11643 => pixel <= "000000";
      when 11644 => pixel <= "000000";
      when 11645 => pixel <= "000000";
      when 11646 => pixel <= "000000";
      when 11647 => pixel <= "000000";
      when 11648 => pixel <= "000000";
      when 11649 => pixel <= "000000";
      when 11650 => pixel <= "000000";
      when 11651 => pixel <= "000000";
      when 11652 => pixel <= "000000";
      when 11653 => pixel <= "000000";
      when 11654 => pixel <= "000000";
      when 11655 => pixel <= "000000";
      when 11656 => pixel <= "000000";
      when 11657 => pixel <= "000000";
      when 11658 => pixel <= "000000";
      when 11659 => pixel <= "000000";
      when 11660 => pixel <= "000000";
      when 11661 => pixel <= "000000";
      when 11662 => pixel <= "000000";
      when 11663 => pixel <= "000000";
      when 11664 => pixel <= "000000";
      when 11665 => pixel <= "000000";
      when 11666 => pixel <= "000000";
      when 11667 => pixel <= "000000";
      when 11668 => pixel <= "000000";
      when 11669 => pixel <= "000000";
      when 11670 => pixel <= "000000";
      when 11671 => pixel <= "000000";
      when 11672 => pixel <= "000000";
      when 11673 => pixel <= "000000";
      when 11674 => pixel <= "000000";
      when 11675 => pixel <= "000000";
      when 11676 => pixel <= "000000";
      when 11677 => pixel <= "000000";
      when 11678 => pixel <= "000000";
      when 11679 => pixel <= "000000";
      when 11680 => pixel <= "000000";
      when 11681 => pixel <= "000000";
      when 11682 => pixel <= "000000";
      when 11683 => pixel <= "000000";
      when 11684 => pixel <= "000000";
      when 11685 => pixel <= "000000";
      when 11686 => pixel <= "000000";
      when 11687 => pixel <= "000000";
      when 11688 => pixel <= "000000";
      when 11689 => pixel <= "000000";
      when 11690 => pixel <= "000000";
      when 11691 => pixel <= "000000";
      when 11692 => pixel <= "000000";
      when 11693 => pixel <= "000000";
      when 11694 => pixel <= "000000";
      when 11695 => pixel <= "000000";
      when 11696 => pixel <= "000000";
      when 11697 => pixel <= "000000";
      when 11698 => pixel <= "000000";
      when 11699 => pixel <= "000000";
      when 11700 => pixel <= "000000";
      when 11701 => pixel <= "000000";
      when 11702 => pixel <= "000000";
      when 11703 => pixel <= "000000";
      when 11704 => pixel <= "000000";
      when 11705 => pixel <= "000000";
      when 11706 => pixel <= "000000";
      when 11707 => pixel <= "000000";
      when 11708 => pixel <= "000000";
      when 11709 => pixel <= "000000";
      when 11710 => pixel <= "000000";
      when 11711 => pixel <= "000000";
      when 11712 => pixel <= "000000";
      when 11713 => pixel <= "000000";
      when 11714 => pixel <= "000000";
      when 11715 => pixel <= "000000";
      when 11716 => pixel <= "000000";
      when 11717 => pixel <= "000000";
      when 11718 => pixel <= "000000";
      when 11719 => pixel <= "000000";
      when 11720 => pixel <= "000000";
      when 11721 => pixel <= "000000";
      when 11722 => pixel <= "000000";
      when 11723 => pixel <= "000000";
      when 11724 => pixel <= "000000";
      when 11725 => pixel <= "000000";
      when 11726 => pixel <= "000000";
      when 11727 => pixel <= "000000";
      when 11728 => pixel <= "000000";
      when 11729 => pixel <= "000000";
      when 11730 => pixel <= "000000";
      when 11731 => pixel <= "000000";
      when 11732 => pixel <= "000000";
      when 11733 => pixel <= "000000";
      when 11734 => pixel <= "000000";
      when 11735 => pixel <= "000000";
      when 11736 => pixel <= "000000";
      when 11737 => pixel <= "000000";
      when 11738 => pixel <= "000000";
      when 11739 => pixel <= "000000";
      when 11740 => pixel <= "000000";
      when 11741 => pixel <= "000000";
      when 11742 => pixel <= "000000";
      when 11743 => pixel <= "000000";
      when 11744 => pixel <= "000000";
      when 11745 => pixel <= "000000";
      when 11746 => pixel <= "000000";
      when 11747 => pixel <= "000000";
      when 11748 => pixel <= "000000";
      when 11749 => pixel <= "000000";
      when 11750 => pixel <= "000000";
      when 11751 => pixel <= "000000";
      when 11752 => pixel <= "000000";
      when 11753 => pixel <= "000000";
      when 11754 => pixel <= "000000";
      when 11755 => pixel <= "000000";
      when 11756 => pixel <= "000000";
      when 11757 => pixel <= "000000";
      when 11758 => pixel <= "000000";
      when 11759 => pixel <= "000000";
      when 11760 => pixel <= "000000";
      when 11761 => pixel <= "000000";
      when 11762 => pixel <= "000000";
      when 11763 => pixel <= "000000";
      when 11764 => pixel <= "000000";
      when 11765 => pixel <= "000000";
      when 11766 => pixel <= "000000";
      when 11767 => pixel <= "000000";
      when 11768 => pixel <= "000000";
      when 11769 => pixel <= "000000";
      when 11770 => pixel <= "000000";
      when 11771 => pixel <= "000000";
      when 11772 => pixel <= "000000";
      when 11773 => pixel <= "000000";
      when 11774 => pixel <= "000000";
      when 11775 => pixel <= "000000";
      when 11776 => pixel <= "000000";
      when 11777 => pixel <= "000000";
      when 11778 => pixel <= "000000";
      when 11779 => pixel <= "000000";
      when 11780 => pixel <= "000000";
      when 11781 => pixel <= "000000";
      when 11782 => pixel <= "000000";
      when 11783 => pixel <= "000000";
      when 11784 => pixel <= "000000";
      when 11785 => pixel <= "000000";
      when 11786 => pixel <= "000000";
      when 11787 => pixel <= "000000";
      when 11788 => pixel <= "000000";
      when 11789 => pixel <= "000000";
      when 11790 => pixel <= "000000";
      when 11791 => pixel <= "000000";
      when 11792 => pixel <= "000000";
      when 11793 => pixel <= "000000";
      when 11794 => pixel <= "000000";
      when 11795 => pixel <= "000000";
      when 11796 => pixel <= "000000";
      when 11797 => pixel <= "000000";
      when 11798 => pixel <= "000000";
      when 11799 => pixel <= "000000";
      when 11800 => pixel <= "000000";
      when 11801 => pixel <= "000000";
      when 11802 => pixel <= "000000";
      when 11803 => pixel <= "000000";
      when 11804 => pixel <= "000000";
      when 11805 => pixel <= "000000";
      when 11806 => pixel <= "000000";
      when 11807 => pixel <= "000000";
      when 11808 => pixel <= "000000";
      when 11809 => pixel <= "000000";
      when 11810 => pixel <= "000000";
      when 11811 => pixel <= "000000";
      when 11812 => pixel <= "000000";
      when 11813 => pixel <= "000000";
      when 11814 => pixel <= "000000";
      when 11815 => pixel <= "000000";
      when 11816 => pixel <= "000000";
      when 11817 => pixel <= "000000";
      when 11818 => pixel <= "000000";
      when 11819 => pixel <= "000000";
      when 11820 => pixel <= "000000";
      when 11821 => pixel <= "000000";
      when 11822 => pixel <= "000000";
      when 11823 => pixel <= "000000";
      when 11824 => pixel <= "000000";
      when 11825 => pixel <= "000000";
      when 11826 => pixel <= "000000";
      when 11827 => pixel <= "000000";
      when 11828 => pixel <= "000000";
      when 11829 => pixel <= "000000";
      when 11830 => pixel <= "000000";
      when 11831 => pixel <= "000000";
      when 11832 => pixel <= "000000";
      when 11833 => pixel <= "000000";
      when 11834 => pixel <= "000000";
      when 11835 => pixel <= "000000";
      when 11836 => pixel <= "000000";
      when 11837 => pixel <= "000000";
      when 11838 => pixel <= "000000";
      when 11839 => pixel <= "000000";
      when 11840 => pixel <= "000000";
      when 11841 => pixel <= "000000";
      when 11842 => pixel <= "000000";
      when 11843 => pixel <= "000000";
      when 11844 => pixel <= "000000";
      when 11845 => pixel <= "000000";
      when 11846 => pixel <= "000000";
      when 11847 => pixel <= "000000";
      when 11848 => pixel <= "000000";
      when 11849 => pixel <= "000000";
      when 11850 => pixel <= "000000";
      when 11851 => pixel <= "000000";
      when 11852 => pixel <= "000000";
      when 11853 => pixel <= "000000";
      when 11854 => pixel <= "000000";
      when 11855 => pixel <= "000000";
      when 11856 => pixel <= "000000";
      when 11857 => pixel <= "000000";
      when 11858 => pixel <= "000000";
      when 11859 => pixel <= "000000";
      when 11860 => pixel <= "000000";
      when 11861 => pixel <= "000000";
      when 11862 => pixel <= "000000";
      when 11863 => pixel <= "000000";
      when 11864 => pixel <= "000000";
      when 11865 => pixel <= "000000";
      when 11866 => pixel <= "000000";
      when 11867 => pixel <= "000000";
      when 11868 => pixel <= "000000";
      when 11869 => pixel <= "000000";
      when 11870 => pixel <= "000000";
      when 11871 => pixel <= "000000";
      when 11872 => pixel <= "000000";
      when 11873 => pixel <= "000000";
      when 11874 => pixel <= "000000";
      when 11875 => pixel <= "000000";
      when 11876 => pixel <= "000000";
      when 11877 => pixel <= "000000";
      when 11878 => pixel <= "000000";
      when 11879 => pixel <= "000000";
      when 11880 => pixel <= "000000";
      when 11881 => pixel <= "000000";
      when 11882 => pixel <= "000000";
      when 11883 => pixel <= "000000";
      when 11884 => pixel <= "000000";
      when 11885 => pixel <= "000000";
      when 11886 => pixel <= "000000";
      when 11887 => pixel <= "000000";
      when 11888 => pixel <= "000000";
      when 11889 => pixel <= "000000";
      when 11890 => pixel <= "000000";
      when 11891 => pixel <= "000000";
      when 11892 => pixel <= "000000";
      when 11893 => pixel <= "000000";
      when 11894 => pixel <= "000000";
      when 11895 => pixel <= "000000";
      when 11896 => pixel <= "000000";
      when 11897 => pixel <= "000000";
      when 11898 => pixel <= "000000";
      when 11899 => pixel <= "000000";
      when 11900 => pixel <= "000000";
      when 11901 => pixel <= "000000";
      when 11902 => pixel <= "000000";
      when 11903 => pixel <= "000000";
      when 11904 => pixel <= "000000";
      when 11905 => pixel <= "000000";
      when 11906 => pixel <= "000000";
      when 11907 => pixel <= "000000";
      when 11908 => pixel <= "000000";
      when 11909 => pixel <= "000000";
      when 11910 => pixel <= "000000";
      when 11911 => pixel <= "000000";
      when 11912 => pixel <= "000000";
      when 11913 => pixel <= "000000";
      when 11914 => pixel <= "000000";
      when 11915 => pixel <= "000000";
      when 11916 => pixel <= "000000";
      when 11917 => pixel <= "000000";
      when 11918 => pixel <= "000000";
      when 11919 => pixel <= "000000";
      when 11920 => pixel <= "000000";
      when 11921 => pixel <= "000000";
      when 11922 => pixel <= "000000";
      when 11923 => pixel <= "000000";
      when 11924 => pixel <= "000000";
      when 11925 => pixel <= "000000";
      when 11926 => pixel <= "000000";
      when 11927 => pixel <= "000000";
      when 11928 => pixel <= "000000";
      when 11929 => pixel <= "000000";
      when 11930 => pixel <= "000000";
      when 11931 => pixel <= "000000";
      when 11932 => pixel <= "000000";
      when 11933 => pixel <= "000000";
      when 11934 => pixel <= "000000";
      when 11935 => pixel <= "000000";
      when 11936 => pixel <= "000000";
      when 11937 => pixel <= "000000";
      when 11938 => pixel <= "000000";
      when 11939 => pixel <= "000000";
      when 11940 => pixel <= "000000";
      when 11941 => pixel <= "000000";
      when 11942 => pixel <= "000000";
      when 11943 => pixel <= "000000";
      when 11944 => pixel <= "000000";
      when 11945 => pixel <= "000000";
      when 11946 => pixel <= "000000";
      when 11947 => pixel <= "000000";
      when 11948 => pixel <= "000000";
      when 11949 => pixel <= "000000";
      when 11950 => pixel <= "000000";
      when 11951 => pixel <= "000000";
      when 11952 => pixel <= "000000";
      when 11953 => pixel <= "000000";
      when 11954 => pixel <= "000000";
      when 11955 => pixel <= "000000";
      when 11956 => pixel <= "000000";
      when 11957 => pixel <= "000000";
      when 11958 => pixel <= "000000";
      when 11959 => pixel <= "000000";
      when 11960 => pixel <= "000000";
      when 11961 => pixel <= "000000";
      when 11962 => pixel <= "000000";
      when 11963 => pixel <= "000000";
      when 11964 => pixel <= "000000";
      when 11965 => pixel <= "000000";
      when 11966 => pixel <= "000000";
      when 11967 => pixel <= "000000";
      when 11968 => pixel <= "000000";
      when 11969 => pixel <= "000000";
      when 11970 => pixel <= "000000";
      when 11971 => pixel <= "000000";
      when 11972 => pixel <= "000000";
      when 11973 => pixel <= "000000";
      when 11974 => pixel <= "000000";
      when 11975 => pixel <= "000000";
      when 11976 => pixel <= "000000";
      when 11977 => pixel <= "000000";
      when 11978 => pixel <= "000000";
      when 11979 => pixel <= "000000";
      when 11980 => pixel <= "000000";
      when 11981 => pixel <= "000000";
      when 11982 => pixel <= "000000";
      when 11983 => pixel <= "000000";
      when 11984 => pixel <= "000000";
      when 11985 => pixel <= "000000";
      when 11986 => pixel <= "000000";
      when 11987 => pixel <= "000000";
      when 11988 => pixel <= "000000";
      when 11989 => pixel <= "000000";
      when 11990 => pixel <= "000000";
      when 11991 => pixel <= "000000";
      when 11992 => pixel <= "000000";
      when 11993 => pixel <= "000000";
      when 11994 => pixel <= "000000";
      when 11995 => pixel <= "000000";
      when 11996 => pixel <= "000000";
      when 11997 => pixel <= "000000";
      when 11998 => pixel <= "000000";
      when 11999 => pixel <= "000000";
      when 12000 => pixel <= "000000";
      when 12001 => pixel <= "000000";
      when 12002 => pixel <= "000000";
      when 12003 => pixel <= "000000";
      when 12004 => pixel <= "000000";
      when 12005 => pixel <= "000000";
      when 12006 => pixel <= "000000";
      when 12007 => pixel <= "000000";
      when 12008 => pixel <= "000000";
      when 12009 => pixel <= "000000";
      when 12010 => pixel <= "000000";
      when 12011 => pixel <= "000000";
      when 12012 => pixel <= "000000";
      when 12013 => pixel <= "000000";
      when 12014 => pixel <= "000000";
      when 12015 => pixel <= "000000";
      when 12016 => pixel <= "000000";
      when 12017 => pixel <= "000000";
      when 12018 => pixel <= "000000";
      when 12019 => pixel <= "000000";
      when 12020 => pixel <= "000000";
      when 12021 => pixel <= "000000";
      when 12022 => pixel <= "000000";
      when 12023 => pixel <= "000000";
      when 12024 => pixel <= "000000";
      when 12025 => pixel <= "000000";
      when 12026 => pixel <= "000000";
      when 12027 => pixel <= "000000";
      when 12028 => pixel <= "000000";
      when 12029 => pixel <= "000000";
      when 12030 => pixel <= "000000";
      when 12031 => pixel <= "000000";
      when 12032 => pixel <= "000000";
      when 12033 => pixel <= "000000";
      when 12034 => pixel <= "000000";
      when 12035 => pixel <= "000000";
      when 12036 => pixel <= "000000";
      when 12037 => pixel <= "000000";
      when 12038 => pixel <= "000000";
      when 12039 => pixel <= "000000";
      when 12040 => pixel <= "000000";
      when 12041 => pixel <= "000000";
      when 12042 => pixel <= "000000";
      when 12043 => pixel <= "000000";
      when 12044 => pixel <= "000000";
      when 12045 => pixel <= "000000";
      when 12046 => pixel <= "000000";
      when 12047 => pixel <= "000000";
      when 12048 => pixel <= "000000";
      when 12049 => pixel <= "000000";
      when 12050 => pixel <= "000000";
      when 12051 => pixel <= "000000";
      when 12052 => pixel <= "000000";
      when 12053 => pixel <= "000000";
      when 12054 => pixel <= "000000";
      when 12055 => pixel <= "000000";
      when 12056 => pixel <= "000000";
      when 12057 => pixel <= "000000";
      when 12058 => pixel <= "000000";
      when 12059 => pixel <= "000000";
      when 12060 => pixel <= "000000";
      when 12061 => pixel <= "000000";
      when 12062 => pixel <= "000000";
      when 12063 => pixel <= "000000";
      when 12064 => pixel <= "000000";
      when 12065 => pixel <= "000000";
      when 12066 => pixel <= "000000";
      when 12067 => pixel <= "000000";
      when 12068 => pixel <= "000000";
      when 12069 => pixel <= "000000";
      when 12070 => pixel <= "000000";
      when 12071 => pixel <= "000000";
      when 12072 => pixel <= "000000";
      when 12073 => pixel <= "000000";
      when 12074 => pixel <= "000000";
      when 12075 => pixel <= "000000";
      when 12076 => pixel <= "000000";
      when 12077 => pixel <= "000000";
      when 12078 => pixel <= "000000";
      when 12079 => pixel <= "000000";
      when 12080 => pixel <= "000000";
      when 12081 => pixel <= "000000";
      when 12082 => pixel <= "000000";
      when 12083 => pixel <= "000000";
      when 12084 => pixel <= "000000";
      when 12085 => pixel <= "000000";
      when 12086 => pixel <= "000000";
      when 12087 => pixel <= "000000";
      when 12088 => pixel <= "000000";
      when 12089 => pixel <= "000000";
      when 12090 => pixel <= "000000";
      when 12091 => pixel <= "000000";
      when 12092 => pixel <= "000000";
      when 12093 => pixel <= "000000";
      when 12094 => pixel <= "000000";
      when 12095 => pixel <= "000000";
      when 12096 => pixel <= "000000";
      when 12097 => pixel <= "000000";
      when 12098 => pixel <= "000000";
      when 12099 => pixel <= "000000";
      when 12100 => pixel <= "000000";
      when 12101 => pixel <= "000000";
      when 12102 => pixel <= "000000";
      when 12103 => pixel <= "000000";
      when 12104 => pixel <= "000000";
      when 12105 => pixel <= "000000";
      when 12106 => pixel <= "000000";
      when 12107 => pixel <= "000000";
      when 12108 => pixel <= "000000";
      when 12109 => pixel <= "000000";
      when 12110 => pixel <= "000000";
      when 12111 => pixel <= "000000";
      when 12112 => pixel <= "000000";
      when 12113 => pixel <= "000000";
      when 12114 => pixel <= "000000";
      when 12115 => pixel <= "000000";
      when 12116 => pixel <= "000000";
      when 12117 => pixel <= "000000";
      when 12118 => pixel <= "000000";
      when 12119 => pixel <= "000000";
      when 12120 => pixel <= "000000";
      when 12121 => pixel <= "000000";
      when 12122 => pixel <= "000000";
      when 12123 => pixel <= "000000";
      when 12124 => pixel <= "000000";
      when 12125 => pixel <= "000000";
      when 12126 => pixel <= "000000";
      when 12127 => pixel <= "000000";
      when 12128 => pixel <= "000000";
      when 12129 => pixel <= "000000";
      when 12130 => pixel <= "000000";
      when 12131 => pixel <= "000000";
      when 12132 => pixel <= "000000";
      when 12133 => pixel <= "000000";
      when 12134 => pixel <= "000000";
      when 12135 => pixel <= "000000";
      when 12136 => pixel <= "000000";
      when 12137 => pixel <= "000000";
      when 12138 => pixel <= "000000";
      when 12139 => pixel <= "000000";
      when 12140 => pixel <= "000000";
      when 12141 => pixel <= "000000";
      when 12142 => pixel <= "000000";
      when 12143 => pixel <= "000000";
      when 12144 => pixel <= "000000";
      when 12145 => pixel <= "000000";
      when 12146 => pixel <= "000000";
      when 12147 => pixel <= "000000";
      when 12148 => pixel <= "000000";
      when 12149 => pixel <= "000000";
      when 12150 => pixel <= "000000";
      when 12151 => pixel <= "000000";
      when 12152 => pixel <= "000000";
      when 12153 => pixel <= "000000";
      when 12154 => pixel <= "000000";
      when 12155 => pixel <= "000000";
      when 12156 => pixel <= "000000";
      when 12157 => pixel <= "000000";
      when 12158 => pixel <= "000000";
      when 12159 => pixel <= "000000";
      when 12160 => pixel <= "000000";
      when 12161 => pixel <= "000000";
      when 12162 => pixel <= "000000";
      when 12163 => pixel <= "000000";
      when 12164 => pixel <= "000000";
      when 12165 => pixel <= "000000";
      when 12166 => pixel <= "000000";
      when 12167 => pixel <= "000000";
      when 12168 => pixel <= "000000";
      when 12169 => pixel <= "000000";
      when 12170 => pixel <= "000000";
      when 12171 => pixel <= "000000";
      when 12172 => pixel <= "000000";
      when 12173 => pixel <= "000000";
      when 12174 => pixel <= "000000";
      when 12175 => pixel <= "000000";
      when 12176 => pixel <= "000000";
      when 12177 => pixel <= "000000";
      when 12178 => pixel <= "000000";
      when 12179 => pixel <= "000000";
      when 12180 => pixel <= "000000";
      when 12181 => pixel <= "000000";
      when 12182 => pixel <= "000000";
      when 12183 => pixel <= "000000";
      when 12184 => pixel <= "000000";
      when 12185 => pixel <= "000000";
      when 12186 => pixel <= "000000";
      when 12187 => pixel <= "000000";
      when 12188 => pixel <= "000000";
      when 12189 => pixel <= "000000";
      when 12190 => pixel <= "000000";
      when 12191 => pixel <= "000000";
      when 12192 => pixel <= "000000";
      when 12193 => pixel <= "000000";
      when 12194 => pixel <= "000000";
      when 12195 => pixel <= "000000";
      when 12196 => pixel <= "000000";
      when 12197 => pixel <= "000000";
      when 12198 => pixel <= "000000";
      when 12199 => pixel <= "000000";
      when 12200 => pixel <= "000000";
      when 12201 => pixel <= "000000";
      when 12202 => pixel <= "000000";
      when 12203 => pixel <= "000000";
      when 12204 => pixel <= "000000";
      when 12205 => pixel <= "000000";
      when 12206 => pixel <= "000000";
      when 12207 => pixel <= "000000";
      when 12208 => pixel <= "000000";
      when 12209 => pixel <= "000000";
      when 12210 => pixel <= "000000";
      when 12211 => pixel <= "000000";
      when 12212 => pixel <= "000000";
      when 12213 => pixel <= "000000";
      when 12214 => pixel <= "000000";
      when 12215 => pixel <= "000000";
      when 12216 => pixel <= "000000";
      when 12217 => pixel <= "000000";
      when 12218 => pixel <= "000000";
      when 12219 => pixel <= "000000";
      when 12220 => pixel <= "000000";
      when 12221 => pixel <= "000000";
      when 12222 => pixel <= "000000";
      when 12223 => pixel <= "000000";
      when 12224 => pixel <= "000000";
      when 12225 => pixel <= "000000";
      when 12226 => pixel <= "000000";
      when 12227 => pixel <= "000000";
      when 12228 => pixel <= "000000";
      when 12229 => pixel <= "000000";
      when 12230 => pixel <= "000000";
      when 12231 => pixel <= "000000";
      when 12232 => pixel <= "000000";
      when 12233 => pixel <= "000000";
      when 12234 => pixel <= "000000";
      when 12235 => pixel <= "000000";
      when 12236 => pixel <= "000000";
      when 12237 => pixel <= "000000";
      when 12238 => pixel <= "000000";
      when 12239 => pixel <= "000000";
      when 12240 => pixel <= "000000";
      when 12241 => pixel <= "000000";
      when 12242 => pixel <= "000000";
      when 12243 => pixel <= "000000";
      when 12244 => pixel <= "000000";
      when 12245 => pixel <= "000000";
      when 12246 => pixel <= "000000";
      when 12247 => pixel <= "000000";
      when 12248 => pixel <= "000000";
      when 12249 => pixel <= "000000";
      when 12250 => pixel <= "000000";
      when 12251 => pixel <= "000000";
      when 12252 => pixel <= "000000";
      when 12253 => pixel <= "000000";
      when 12254 => pixel <= "000000";
      when 12255 => pixel <= "000000";
      when 12256 => pixel <= "000000";
      when 12257 => pixel <= "000000";
      when 12258 => pixel <= "000000";
      when 12259 => pixel <= "000000";
      when 12260 => pixel <= "000000";
      when 12261 => pixel <= "000000";
      when 12262 => pixel <= "000000";
      when 12263 => pixel <= "000000";
      when 12264 => pixel <= "000000";
      when 12265 => pixel <= "000000";
      when 12266 => pixel <= "000000";
      when 12267 => pixel <= "000000";
      when 12268 => pixel <= "000000";
      when 12269 => pixel <= "000000";
      when 12270 => pixel <= "000000";
      when 12271 => pixel <= "000000";
      when 12272 => pixel <= "000000";
      when 12273 => pixel <= "000000";
      when 12274 => pixel <= "000000";
      when 12275 => pixel <= "000000";
      when 12276 => pixel <= "000000";
      when 12277 => pixel <= "000000";
      when 12278 => pixel <= "000000";
      when 12279 => pixel <= "000000";
      when 12280 => pixel <= "000000";
      when 12281 => pixel <= "000000";
      when 12282 => pixel <= "000000";
      when 12283 => pixel <= "000000";
      when 12284 => pixel <= "000000";
      when 12285 => pixel <= "000000";
      when 12286 => pixel <= "000000";
      when 12287 => pixel <= "000000";
      when 12288 => pixel <= "000000";
      when 12289 => pixel <= "000000";
      when 12290 => pixel <= "000000";
      when 12291 => pixel <= "000000";
      when 12292 => pixel <= "000000";
      when 12293 => pixel <= "000000";
      when 12294 => pixel <= "000000";
      when 12295 => pixel <= "000000";
      when 12296 => pixel <= "000000";
      when 12297 => pixel <= "000000";
      when 12298 => pixel <= "000000";
      when 12299 => pixel <= "000000";
      when 12300 => pixel <= "000000";
      when 12301 => pixel <= "000000";
      when 12302 => pixel <= "000000";
      when 12303 => pixel <= "000000";
      when 12304 => pixel <= "000000";
      when 12305 => pixel <= "000000";
      when 12306 => pixel <= "000000";
      when 12307 => pixel <= "000000";
      when 12308 => pixel <= "000000";
      when 12309 => pixel <= "000000";
      when 12310 => pixel <= "000000";
      when 12311 => pixel <= "000000";
      when 12312 => pixel <= "000000";
      when 12313 => pixel <= "000000";
      when 12314 => pixel <= "000000";
      when 12315 => pixel <= "000000";
      when 12316 => pixel <= "000000";
      when 12317 => pixel <= "000000";
      when 12318 => pixel <= "000000";
      when 12319 => pixel <= "000000";
      when 12320 => pixel <= "000000";
      when 12321 => pixel <= "000000";
      when 12322 => pixel <= "000000";
      when 12323 => pixel <= "000000";
      when 12324 => pixel <= "000000";
      when 12325 => pixel <= "000000";
      when 12326 => pixel <= "000000";
      when 12327 => pixel <= "000000";
      when 12328 => pixel <= "000000";
      when 12329 => pixel <= "000000";
      when 12330 => pixel <= "000000";
      when 12331 => pixel <= "000000";
      when 12332 => pixel <= "000000";
      when 12333 => pixel <= "000000";
      when 12334 => pixel <= "000000";
      when 12335 => pixel <= "000000";
      when 12336 => pixel <= "000000";
      when 12337 => pixel <= "000000";
      when 12338 => pixel <= "000000";
      when 12339 => pixel <= "000000";
      when 12340 => pixel <= "000000";
      when 12341 => pixel <= "000000";
      when 12342 => pixel <= "000000";
      when 12343 => pixel <= "000000";
      when 12344 => pixel <= "000000";
      when 12345 => pixel <= "000000";
      when 12346 => pixel <= "000000";
      when 12347 => pixel <= "000000";
      when 12348 => pixel <= "000000";
      when 12349 => pixel <= "000000";
      when 12350 => pixel <= "000000";
      when 12351 => pixel <= "000000";
      when 12352 => pixel <= "000000";
      when 12353 => pixel <= "000000";
      when 12354 => pixel <= "000000";
      when 12355 => pixel <= "000000";
      when 12356 => pixel <= "000000";
      when 12357 => pixel <= "000000";
      when 12358 => pixel <= "000000";
      when 12359 => pixel <= "000000";
      when 12360 => pixel <= "000000";
      when 12361 => pixel <= "000000";
      when 12362 => pixel <= "000000";
      when 12363 => pixel <= "000000";
      when 12364 => pixel <= "000000";
      when 12365 => pixel <= "000000";
      when 12366 => pixel <= "000000";
      when 12367 => pixel <= "000000";
      when 12368 => pixel <= "000000";
      when 12369 => pixel <= "000000";
      when 12370 => pixel <= "000000";
      when 12371 => pixel <= "000000";
      when 12372 => pixel <= "000000";
      when 12373 => pixel <= "000000";
      when 12374 => pixel <= "000000";
      when 12375 => pixel <= "000000";
      when 12376 => pixel <= "000000";
      when 12377 => pixel <= "000000";
      when 12378 => pixel <= "000000";
      when 12379 => pixel <= "000000";
      when 12380 => pixel <= "000000";
      when 12381 => pixel <= "000000";
      when 12382 => pixel <= "000000";
      when 12383 => pixel <= "000000";
      when 12384 => pixel <= "000000";
      when 12385 => pixel <= "000000";
      when 12386 => pixel <= "000000";
      when 12387 => pixel <= "000000";
      when 12388 => pixel <= "000000";
      when 12389 => pixel <= "000000";
      when 12390 => pixel <= "000000";
      when 12391 => pixel <= "000000";
      when 12392 => pixel <= "000000";
      when 12393 => pixel <= "000000";
      when 12394 => pixel <= "000000";
      when 12395 => pixel <= "000000";
      when 12396 => pixel <= "000000";
      when 12397 => pixel <= "000000";
      when 12398 => pixel <= "000000";
      when 12399 => pixel <= "000000";
      when 12400 => pixel <= "000000";
      when 12401 => pixel <= "000000";
      when 12402 => pixel <= "000000";
      when 12403 => pixel <= "000000";
      when 12404 => pixel <= "000000";
      when 12405 => pixel <= "000000";
      when 12406 => pixel <= "000000";
      when 12407 => pixel <= "000000";
      when 12408 => pixel <= "000000";
      when 12409 => pixel <= "000000";
      when 12410 => pixel <= "000000";
      when 12411 => pixel <= "000000";
      when 12412 => pixel <= "000000";
      when 12413 => pixel <= "000000";
      when 12414 => pixel <= "000000";
      when 12415 => pixel <= "000000";
      when 12416 => pixel <= "000000";
      when 12417 => pixel <= "000000";
      when 12418 => pixel <= "000000";
      when 12419 => pixel <= "000000";
      when 12420 => pixel <= "000000";
      when 12421 => pixel <= "000000";
      when 12422 => pixel <= "000000";
      when 12423 => pixel <= "000000";
      when 12424 => pixel <= "000000";
      when 12425 => pixel <= "000000";
      when 12426 => pixel <= "000000";
      when 12427 => pixel <= "000000";
      when 12428 => pixel <= "000000";
      when 12429 => pixel <= "000000";
      when 12430 => pixel <= "000000";
      when 12431 => pixel <= "000000";
      when 12432 => pixel <= "000000";
      when 12433 => pixel <= "000000";
      when 12434 => pixel <= "000000";
      when 12435 => pixel <= "000000";
      when 12436 => pixel <= "000000";
      when 12437 => pixel <= "000000";
      when 12438 => pixel <= "000000";
      when 12439 => pixel <= "000000";
      when 12440 => pixel <= "000000";
      when 12441 => pixel <= "000000";
      when 12442 => pixel <= "000000";
      when 12443 => pixel <= "000000";
      when 12444 => pixel <= "000000";
      when 12445 => pixel <= "000000";
      when 12446 => pixel <= "000000";
      when 12447 => pixel <= "000000";
      when 12448 => pixel <= "000000";
      when 12449 => pixel <= "000000";
      when 12450 => pixel <= "000000";
      when 12451 => pixel <= "000000";
      when 12452 => pixel <= "000000";
      when 12453 => pixel <= "000000";
      when 12454 => pixel <= "000000";
      when 12455 => pixel <= "000000";
      when 12456 => pixel <= "000000";
      when 12457 => pixel <= "000000";
      when 12458 => pixel <= "000000";
      when 12459 => pixel <= "000000";
      when 12460 => pixel <= "000000";
      when 12461 => pixel <= "000000";
      when 12462 => pixel <= "000000";
      when 12463 => pixel <= "000000";
      when 12464 => pixel <= "000000";
      when 12465 => pixel <= "000000";
      when 12466 => pixel <= "000000";
      when 12467 => pixel <= "000000";
      when 12468 => pixel <= "000000";
      when 12469 => pixel <= "000000";
      when 12470 => pixel <= "000000";
      when 12471 => pixel <= "000000";
      when 12472 => pixel <= "000000";
      when 12473 => pixel <= "000000";
      when 12474 => pixel <= "000000";
      when 12475 => pixel <= "000000";
      when 12476 => pixel <= "000000";
      when 12477 => pixel <= "000000";
      when 12478 => pixel <= "000000";
      when 12479 => pixel <= "000000";
      when 12480 => pixel <= "000000";
      when 12481 => pixel <= "000000";
      when 12482 => pixel <= "000000";
      when 12483 => pixel <= "000000";
      when 12484 => pixel <= "000000";
      when 12485 => pixel <= "000000";
      when 12486 => pixel <= "000000";
      when 12487 => pixel <= "000000";
      when 12488 => pixel <= "000000";
      when 12489 => pixel <= "000000";
      when 12490 => pixel <= "000000";
      when 12491 => pixel <= "000000";
      when 12492 => pixel <= "000000";
      when 12493 => pixel <= "000000";
      when 12494 => pixel <= "000000";
      when 12495 => pixel <= "000000";
      when 12496 => pixel <= "000000";
      when 12497 => pixel <= "000000";
      when 12498 => pixel <= "000000";
      when 12499 => pixel <= "000000";
      when 12500 => pixel <= "000000";
      when 12501 => pixel <= "000000";
      when 12502 => pixel <= "000000";
      when 12503 => pixel <= "000000";
      when 12504 => pixel <= "000000";
      when 12505 => pixel <= "000000";
      when 12506 => pixel <= "000000";
      when 12507 => pixel <= "000000";
      when 12508 => pixel <= "000000";
      when 12509 => pixel <= "000000";
      when 12510 => pixel <= "000000";
      when 12511 => pixel <= "000000";
      when 12512 => pixel <= "000000";
      when 12513 => pixel <= "000000";
      when 12514 => pixel <= "000000";
      when 12515 => pixel <= "000000";
      when 12516 => pixel <= "000000";
      when 12517 => pixel <= "000000";
      when 12518 => pixel <= "000000";
      when 12519 => pixel <= "000000";
      when 12520 => pixel <= "000000";
      when 12521 => pixel <= "000000";
      when 12522 => pixel <= "000000";
      when 12523 => pixel <= "000000";
      when 12524 => pixel <= "000000";
      when 12525 => pixel <= "000000";
      when 12526 => pixel <= "000000";
      when 12527 => pixel <= "000000";
      when 12528 => pixel <= "000000";
      when 12529 => pixel <= "000000";
      when 12530 => pixel <= "000000";
      when 12531 => pixel <= "000000";
      when 12532 => pixel <= "000000";
      when 12533 => pixel <= "000000";
      when 12534 => pixel <= "000000";
      when 12535 => pixel <= "000000";
      when 12536 => pixel <= "000000";
      when 12537 => pixel <= "000000";
      when 12538 => pixel <= "000000";
      when 12539 => pixel <= "000000";
      when 12540 => pixel <= "000000";
      when 12541 => pixel <= "000000";
      when 12542 => pixel <= "000000";
      when 12543 => pixel <= "000000";
      when 12544 => pixel <= "000000";
      when 12545 => pixel <= "000000";
      when 12546 => pixel <= "000000";
      when 12547 => pixel <= "000000";
      when 12548 => pixel <= "000000";
      when 12549 => pixel <= "000000";
      when 12550 => pixel <= "000000";
      when 12551 => pixel <= "000000";
      when 12552 => pixel <= "000000";
      when 12553 => pixel <= "000000";
      when 12554 => pixel <= "000000";
      when 12555 => pixel <= "000000";
      when 12556 => pixel <= "000000";
      when 12557 => pixel <= "000000";
      when 12558 => pixel <= "000000";
      when 12559 => pixel <= "000000";
      when 12560 => pixel <= "000000";
      when 12561 => pixel <= "000000";
      when 12562 => pixel <= "000000";
      when 12563 => pixel <= "000000";
      when 12564 => pixel <= "000000";
      when 12565 => pixel <= "000000";
      when 12566 => pixel <= "000000";
      when 12567 => pixel <= "000000";
      when 12568 => pixel <= "000000";
      when 12569 => pixel <= "000000";
      when 12570 => pixel <= "000000";
      when 12571 => pixel <= "000000";
      when 12572 => pixel <= "000000";
      when 12573 => pixel <= "000000";
      when 12574 => pixel <= "000000";
      when 12575 => pixel <= "000000";
      when 12576 => pixel <= "000000";
      when 12577 => pixel <= "000000";
      when 12578 => pixel <= "000000";
      when 12579 => pixel <= "000000";
      when 12580 => pixel <= "000000";
      when 12581 => pixel <= "000000";
      when 12582 => pixel <= "000000";
      when 12583 => pixel <= "000000";
      when 12584 => pixel <= "000000";
      when 12585 => pixel <= "000000";
      when 12586 => pixel <= "000000";
      when 12587 => pixel <= "000000";
      when 12588 => pixel <= "000000";
      when 12589 => pixel <= "000000";
      when 12590 => pixel <= "000000";
      when 12591 => pixel <= "000000";
      when 12592 => pixel <= "000000";
      when 12593 => pixel <= "000000";
      when 12594 => pixel <= "000000";
      when 12595 => pixel <= "000000";
      when 12596 => pixel <= "000000";
      when 12597 => pixel <= "000000";
      when 12598 => pixel <= "000000";
      when 12599 => pixel <= "000000";
      when 12600 => pixel <= "000000";
      when 12601 => pixel <= "000000";
      when 12602 => pixel <= "000000";
      when 12603 => pixel <= "000000";
      when 12604 => pixel <= "000000";
      when 12605 => pixel <= "000000";
      when 12606 => pixel <= "000000";
      when 12607 => pixel <= "000000";
      when 12608 => pixel <= "000000";
      when 12609 => pixel <= "000000";
      when 12610 => pixel <= "000000";
      when 12611 => pixel <= "000000";
      when 12612 => pixel <= "000000";
      when 12613 => pixel <= "000000";
      when 12614 => pixel <= "000000";
      when 12615 => pixel <= "000000";
      when 12616 => pixel <= "000000";
      when 12617 => pixel <= "000000";
      when 12618 => pixel <= "000000";
      when 12619 => pixel <= "000000";
      when 12620 => pixel <= "000000";
      when 12621 => pixel <= "000000";
      when 12622 => pixel <= "000000";
      when 12623 => pixel <= "000000";
      when 12624 => pixel <= "000000";
      when 12625 => pixel <= "000000";
      when 12626 => pixel <= "000000";
      when 12627 => pixel <= "000000";
      when 12628 => pixel <= "000000";
      when 12629 => pixel <= "000000";
      when 12630 => pixel <= "000000";
      when 12631 => pixel <= "000000";
      when 12632 => pixel <= "000000";
      when 12633 => pixel <= "000000";
      when 12634 => pixel <= "000000";
      when 12635 => pixel <= "000000";
      when 12636 => pixel <= "000000";
      when 12637 => pixel <= "000000";
      when 12638 => pixel <= "000000";
      when 12639 => pixel <= "000000";
      when 12640 => pixel <= "000000";
      when 12641 => pixel <= "000000";
      when 12642 => pixel <= "000000";
      when 12643 => pixel <= "000000";
      when 12644 => pixel <= "000000";
      when 12645 => pixel <= "000000";
      when 12646 => pixel <= "000000";
      when 12647 => pixel <= "000000";
      when 12648 => pixel <= "000000";
      when 12649 => pixel <= "000000";
      when 12650 => pixel <= "000000";
      when 12651 => pixel <= "000000";
      when 12652 => pixel <= "000000";
      when 12653 => pixel <= "000000";
      when 12654 => pixel <= "000000";
      when 12655 => pixel <= "000000";
      when 12656 => pixel <= "000000";
      when 12657 => pixel <= "000000";
      when 12658 => pixel <= "000000";
      when 12659 => pixel <= "000000";
      when 12660 => pixel <= "000000";
      when 12661 => pixel <= "000000";
      when 12662 => pixel <= "000000";
      when 12663 => pixel <= "000000";
      when 12664 => pixel <= "000000";
      when 12665 => pixel <= "000000";
      when 12666 => pixel <= "000000";
      when 12667 => pixel <= "000000";
      when 12668 => pixel <= "000000";
      when 12669 => pixel <= "000000";
      when 12670 => pixel <= "000000";
      when 12671 => pixel <= "000000";
      when 12672 => pixel <= "000000";
      when 12673 => pixel <= "000000";
      when 12674 => pixel <= "000000";
      when 12675 => pixel <= "000000";
      when 12676 => pixel <= "000000";
      when 12677 => pixel <= "000000";
      when 12678 => pixel <= "000000";
      when 12679 => pixel <= "000000";
      when 12680 => pixel <= "000000";
      when 12681 => pixel <= "000000";
      when 12682 => pixel <= "000000";
      when 12683 => pixel <= "000000";
      when 12684 => pixel <= "000000";
      when 12685 => pixel <= "000000";
      when 12686 => pixel <= "000000";
      when 12687 => pixel <= "000000";
      when 12688 => pixel <= "000000";
      when 12689 => pixel <= "000000";
      when 12690 => pixel <= "000000";
      when 12691 => pixel <= "000000";
      when 12692 => pixel <= "000000";
      when 12693 => pixel <= "000000";
      when 12694 => pixel <= "000000";
      when 12695 => pixel <= "000000";
      when 12696 => pixel <= "000000";
      when 12697 => pixel <= "000000";
      when 12698 => pixel <= "000000";
      when 12699 => pixel <= "000000";
      when 12700 => pixel <= "000000";
      when 12701 => pixel <= "000000";
      when 12702 => pixel <= "000000";
      when 12703 => pixel <= "000000";
      when 12704 => pixel <= "000000";
      when 12705 => pixel <= "000000";
      when 12706 => pixel <= "000000";
      when 12707 => pixel <= "000000";
      when 12708 => pixel <= "000000";
      when 12709 => pixel <= "000000";
      when 12710 => pixel <= "000000";
      when 12711 => pixel <= "000000";
      when 12712 => pixel <= "000000";
      when 12713 => pixel <= "000000";
      when 12714 => pixel <= "000000";
      when 12715 => pixel <= "000000";
      when 12716 => pixel <= "000000";
      when 12717 => pixel <= "000000";
      when 12718 => pixel <= "000000";
      when 12719 => pixel <= "000000";
      when 12720 => pixel <= "000000";
      when 12721 => pixel <= "000000";
      when 12722 => pixel <= "000000";
      when 12723 => pixel <= "000000";
      when 12724 => pixel <= "000000";
      when 12725 => pixel <= "000000";
      when 12726 => pixel <= "000000";
      when 12727 => pixel <= "000000";
      when 12728 => pixel <= "000000";
      when 12729 => pixel <= "000000";
      when 12730 => pixel <= "000000";
      when 12731 => pixel <= "000000";
      when 12732 => pixel <= "000000";
      when 12733 => pixel <= "000000";
      when 12734 => pixel <= "000000";
      when 12735 => pixel <= "000000";
      when 12736 => pixel <= "000000";
      when 12737 => pixel <= "000000";
      when 12738 => pixel <= "000000";
      when 12739 => pixel <= "000000";
      when 12740 => pixel <= "000000";
      when 12741 => pixel <= "000000";
      when 12742 => pixel <= "000000";
      when 12743 => pixel <= "000000";
      when 12744 => pixel <= "000000";
      when 12745 => pixel <= "000000";
      when 12746 => pixel <= "000000";
      when 12747 => pixel <= "000000";
      when 12748 => pixel <= "000000";
      when 12749 => pixel <= "000000";
      when 12750 => pixel <= "000000";
      when 12751 => pixel <= "000000";
      when 12752 => pixel <= "000000";
      when 12753 => pixel <= "000000";
      when 12754 => pixel <= "000000";
      when 12755 => pixel <= "000000";
      when 12756 => pixel <= "000000";
      when 12757 => pixel <= "000000";
      when 12758 => pixel <= "000000";
      when 12759 => pixel <= "000000";
      when 12760 => pixel <= "000000";
      when 12761 => pixel <= "000000";
      when 12762 => pixel <= "000000";
      when 12763 => pixel <= "000000";
      when 12764 => pixel <= "000000";
      when 12765 => pixel <= "000000";
      when 12766 => pixel <= "000000";
      when 12767 => pixel <= "000000";
      when 12768 => pixel <= "000000";
      when 12769 => pixel <= "000000";
      when 12770 => pixel <= "000000";
      when 12771 => pixel <= "000000";
      when 12772 => pixel <= "000000";
      when 12773 => pixel <= "000000";
      when 12774 => pixel <= "000000";
      when 12775 => pixel <= "000000";
      when 12776 => pixel <= "000000";
      when 12777 => pixel <= "000000";
      when 12778 => pixel <= "000000";
      when 12779 => pixel <= "000000";
      when 12780 => pixel <= "000000";
      when 12781 => pixel <= "000000";
      when 12782 => pixel <= "000000";
      when 12783 => pixel <= "000000";
      when 12784 => pixel <= "000000";
      when 12785 => pixel <= "000000";
      when 12786 => pixel <= "000000";
      when 12787 => pixel <= "000000";
      when 12788 => pixel <= "000000";
      when 12789 => pixel <= "000000";
      when 12790 => pixel <= "000000";
      when 12791 => pixel <= "000000";
      when 12792 => pixel <= "000000";
      when 12793 => pixel <= "000000";
      when 12794 => pixel <= "000000";
      when 12795 => pixel <= "000000";
      when 12796 => pixel <= "000000";
      when 12797 => pixel <= "000000";
      when 12798 => pixel <= "000000";
      when 12799 => pixel <= "000000";
      when 12800 => pixel <= "000000";
      when 12801 => pixel <= "000000";
      when 12802 => pixel <= "000000";
      when 12803 => pixel <= "000000";
      when 12804 => pixel <= "000000";
      when 12805 => pixel <= "000000";
      when 12806 => pixel <= "000000";
      when 12807 => pixel <= "000000";
      when 12808 => pixel <= "000000";
      when 12809 => pixel <= "000000";
      when 12810 => pixel <= "000000";
      when 12811 => pixel <= "000000";
      when 12812 => pixel <= "000000";
      when 12813 => pixel <= "000000";
      when 12814 => pixel <= "000000";
      when 12815 => pixel <= "000000";
      when 12816 => pixel <= "000000";
      when 12817 => pixel <= "000000";
      when 12818 => pixel <= "000000";
      when 12819 => pixel <= "000000";
      when 12820 => pixel <= "000000";
      when 12821 => pixel <= "000000";
      when 12822 => pixel <= "000000";
      when 12823 => pixel <= "000000";
      when 12824 => pixel <= "000000";
      when 12825 => pixel <= "000000";
      when 12826 => pixel <= "000000";
      when 12827 => pixel <= "000000";
      when 12828 => pixel <= "000000";
      when 12829 => pixel <= "000000";
      when 12830 => pixel <= "000000";
      when 12831 => pixel <= "000000";
      when 12832 => pixel <= "000000";
      when 12833 => pixel <= "000000";
      when 12834 => pixel <= "000000";
      when 12835 => pixel <= "000000";
      when 12836 => pixel <= "000000";
      when 12837 => pixel <= "000000";
      when 12838 => pixel <= "000000";
      when 12839 => pixel <= "000000";
      when 12840 => pixel <= "000000";
      when 12841 => pixel <= "000000";
      when 12842 => pixel <= "000000";
      when 12843 => pixel <= "000000";
      when 12844 => pixel <= "000000";
      when 12845 => pixel <= "000000";
      when 12846 => pixel <= "000000";
      when 12847 => pixel <= "000000";
      when 12848 => pixel <= "000000";
      when 12849 => pixel <= "000000";
      when 12850 => pixel <= "000000";
      when 12851 => pixel <= "000000";
      when 12852 => pixel <= "000000";
      when 12853 => pixel <= "000000";
      when 12854 => pixel <= "000000";
      when 12855 => pixel <= "000000";
      when 12856 => pixel <= "000000";
      when 12857 => pixel <= "000000";
      when 12858 => pixel <= "000000";
      when 12859 => pixel <= "000000";
      when 12860 => pixel <= "000000";
      when 12861 => pixel <= "000000";
      when 12862 => pixel <= "000000";
      when 12863 => pixel <= "000000";
      when 12864 => pixel <= "000000";
      when 12865 => pixel <= "000000";
      when 12866 => pixel <= "000000";
      when 12867 => pixel <= "000000";
      when 12868 => pixel <= "000000";
      when 12869 => pixel <= "000000";
      when 12870 => pixel <= "000000";
      when 12871 => pixel <= "000000";
      when 12872 => pixel <= "000000";
      when 12873 => pixel <= "000000";
      when 12874 => pixel <= "000000";
      when 12875 => pixel <= "000000";
      when 12876 => pixel <= "000000";
      when 12877 => pixel <= "000000";
      when 12878 => pixel <= "000000";
      when 12879 => pixel <= "000000";
      when 12880 => pixel <= "000000";
      when 12881 => pixel <= "000000";
      when 12882 => pixel <= "000000";
      when 12883 => pixel <= "000000";
      when 12884 => pixel <= "000000";
      when 12885 => pixel <= "000000";
      when 12886 => pixel <= "000000";
      when 12887 => pixel <= "000000";
      when 12888 => pixel <= "000000";
      when 12889 => pixel <= "000000";
      when 12890 => pixel <= "000000";
      when 12891 => pixel <= "000000";
      when 12892 => pixel <= "000000";
      when 12893 => pixel <= "000000";
      when 12894 => pixel <= "000000";
      when 12895 => pixel <= "000000";
      when 12896 => pixel <= "000000";
      when 12897 => pixel <= "000000";
      when 12898 => pixel <= "000000";
      when 12899 => pixel <= "000000";
      when 12900 => pixel <= "000000";
      when 12901 => pixel <= "000000";
      when 12902 => pixel <= "000000";
      when 12903 => pixel <= "000000";
      when 12904 => pixel <= "000000";
      when 12905 => pixel <= "000000";
      when 12906 => pixel <= "000000";
      when 12907 => pixel <= "000000";
      when 12908 => pixel <= "000000";
      when 12909 => pixel <= "000000";
      when 12910 => pixel <= "000000";
      when 12911 => pixel <= "000000";
      when 12912 => pixel <= "000000";
      when 12913 => pixel <= "000000";
      when 12914 => pixel <= "000000";
      when 12915 => pixel <= "000000";
      when 12916 => pixel <= "000000";
      when 12917 => pixel <= "000000";
      when 12918 => pixel <= "000000";
      when 12919 => pixel <= "000000";
      when 12920 => pixel <= "000000";
      when 12921 => pixel <= "000000";
      when 12922 => pixel <= "000000";
      when 12923 => pixel <= "000000";
      when 12924 => pixel <= "000000";
      when 12925 => pixel <= "000000";
      when 12926 => pixel <= "000000";
      when 12927 => pixel <= "000000";
      when 12928 => pixel <= "000000";
      when 12929 => pixel <= "000000";
      when 12930 => pixel <= "000000";
      when 12931 => pixel <= "000000";
      when 12932 => pixel <= "000000";
      when 12933 => pixel <= "000000";
      when 12934 => pixel <= "000000";
      when 12935 => pixel <= "000000";
      when 12936 => pixel <= "000000";
      when 12937 => pixel <= "000000";
      when 12938 => pixel <= "000000";
      when 12939 => pixel <= "000000";
      when 12940 => pixel <= "000000";
      when 12941 => pixel <= "000000";
      when 12942 => pixel <= "000000";
      when 12943 => pixel <= "000000";
      when 12944 => pixel <= "000000";
      when 12945 => pixel <= "000000";
      when 12946 => pixel <= "000000";
      when 12947 => pixel <= "000000";
      when 12948 => pixel <= "000000";
      when 12949 => pixel <= "000000";
      when 12950 => pixel <= "000000";
      when 12951 => pixel <= "000000";
      when 12952 => pixel <= "000000";
      when 12953 => pixel <= "000000";
      when 12954 => pixel <= "000000";
      when 12955 => pixel <= "000000";
      when 12956 => pixel <= "000000";
      when 12957 => pixel <= "000000";
      when 12958 => pixel <= "000000";
      when 12959 => pixel <= "000000";
      when 12960 => pixel <= "000000";
      when 12961 => pixel <= "000000";
      when 12962 => pixel <= "000000";
      when 12963 => pixel <= "000000";
      when 12964 => pixel <= "000000";
      when 12965 => pixel <= "000000";
      when 12966 => pixel <= "000000";
      when 12967 => pixel <= "000000";
      when 12968 => pixel <= "000000";
      when 12969 => pixel <= "000000";
      when 12970 => pixel <= "000000";
      when 12971 => pixel <= "000000";
      when 12972 => pixel <= "000000";
      when 12973 => pixel <= "000000";
      when 12974 => pixel <= "000000";
      when 12975 => pixel <= "000000";
      when 12976 => pixel <= "000000";
      when 12977 => pixel <= "000000";
      when 12978 => pixel <= "000000";
      when 12979 => pixel <= "000000";
      when 12980 => pixel <= "000000";
      when 12981 => pixel <= "000000";
      when 12982 => pixel <= "000000";
      when 12983 => pixel <= "000000";
      when 12984 => pixel <= "000000";
      when 12985 => pixel <= "000000";
      when 12986 => pixel <= "000000";
      when 12987 => pixel <= "000000";
      when 12988 => pixel <= "000000";
      when 12989 => pixel <= "000000";
      when 12990 => pixel <= "000000";
      when 12991 => pixel <= "000000";
      when 12992 => pixel <= "000000";
      when 12993 => pixel <= "000000";
      when 12994 => pixel <= "000000";
      when 12995 => pixel <= "000000";
      when 12996 => pixel <= "000000";
      when 12997 => pixel <= "000000";
      when 12998 => pixel <= "000000";
      when 12999 => pixel <= "000000";
      when 13000 => pixel <= "000000";
      when 13001 => pixel <= "000000";
      when 13002 => pixel <= "000000";
      when 13003 => pixel <= "000000";
      when 13004 => pixel <= "000000";
      when 13005 => pixel <= "000000";
      when 13006 => pixel <= "000000";
      when 13007 => pixel <= "000000";
      when 13008 => pixel <= "000000";
      when 13009 => pixel <= "000000";
      when 13010 => pixel <= "000000";
      when 13011 => pixel <= "000000";
      when 13012 => pixel <= "000000";
      when 13013 => pixel <= "000000";
      when 13014 => pixel <= "000000";
      when 13015 => pixel <= "000000";
      when 13016 => pixel <= "000000";
      when 13017 => pixel <= "000000";
      when 13018 => pixel <= "000000";
      when 13019 => pixel <= "000000";
      when 13020 => pixel <= "000000";
      when 13021 => pixel <= "000000";
      when 13022 => pixel <= "000000";
      when 13023 => pixel <= "000000";
      when 13024 => pixel <= "000000";
      when 13025 => pixel <= "000000";
      when 13026 => pixel <= "000000";
      when 13027 => pixel <= "000000";
      when 13028 => pixel <= "000000";
      when 13029 => pixel <= "000000";
      when 13030 => pixel <= "000000";
      when 13031 => pixel <= "000000";
      when 13032 => pixel <= "000000";
      when 13033 => pixel <= "000000";
      when 13034 => pixel <= "000000";
      when 13035 => pixel <= "000000";
      when 13036 => pixel <= "000000";
      when 13037 => pixel <= "000000";
      when 13038 => pixel <= "000000";
      when 13039 => pixel <= "000000";
      when 13040 => pixel <= "000000";
      when 13041 => pixel <= "000000";
      when 13042 => pixel <= "000000";
      when 13043 => pixel <= "000000";
      when 13044 => pixel <= "000000";
      when 13045 => pixel <= "000000";
      when 13046 => pixel <= "000000";
      when 13047 => pixel <= "000000";
      when 13048 => pixel <= "000000";
      when 13049 => pixel <= "000000";
      when 13050 => pixel <= "000000";
      when 13051 => pixel <= "000000";
      when 13052 => pixel <= "000000";
      when 13053 => pixel <= "000000";
      when 13054 => pixel <= "000000";
      when 13055 => pixel <= "000000";
      when 13056 => pixel <= "000000";
      when 13057 => pixel <= "000000";
      when 13058 => pixel <= "000000";
      when 13059 => pixel <= "000000";
      when 13060 => pixel <= "000000";
      when 13061 => pixel <= "000000";
      when 13062 => pixel <= "000000";
      when 13063 => pixel <= "000000";
      when 13064 => pixel <= "000000";
      when 13065 => pixel <= "000000";
      when 13066 => pixel <= "000000";
      when 13067 => pixel <= "000000";
      when 13068 => pixel <= "000000";
      when 13069 => pixel <= "000000";
      when 13070 => pixel <= "000000";
      when 13071 => pixel <= "000000";
      when 13072 => pixel <= "000000";
      when 13073 => pixel <= "000000";
      when 13074 => pixel <= "000000";
      when 13075 => pixel <= "000000";
      when 13076 => pixel <= "000000";
      when 13077 => pixel <= "000000";
      when 13078 => pixel <= "000000";
      when 13079 => pixel <= "000000";
      when 13080 => pixel <= "000000";
      when 13081 => pixel <= "000000";
      when 13082 => pixel <= "000000";
      when 13083 => pixel <= "000000";
      when 13084 => pixel <= "000000";
      when 13085 => pixel <= "000000";
      when 13086 => pixel <= "000000";
      when 13087 => pixel <= "000000";
      when 13088 => pixel <= "000000";
      when 13089 => pixel <= "000000";
      when 13090 => pixel <= "000000";
      when 13091 => pixel <= "000000";
      when 13092 => pixel <= "000000";
      when 13093 => pixel <= "000000";
      when 13094 => pixel <= "000000";
      when 13095 => pixel <= "000000";
      when 13096 => pixel <= "000000";
      when 13097 => pixel <= "000000";
      when 13098 => pixel <= "000000";
      when 13099 => pixel <= "000000";
      when 13100 => pixel <= "000000";
      when 13101 => pixel <= "000000";
      when 13102 => pixel <= "000000";
      when 13103 => pixel <= "000000";
      when 13104 => pixel <= "000000";
      when 13105 => pixel <= "000000";
      when 13106 => pixel <= "000000";
      when 13107 => pixel <= "000000";
      when 13108 => pixel <= "000000";
      when 13109 => pixel <= "000000";
      when 13110 => pixel <= "000000";
      when 13111 => pixel <= "000000";
      when 13112 => pixel <= "000000";
      when 13113 => pixel <= "000000";
      when 13114 => pixel <= "000000";
      when 13115 => pixel <= "000000";
      when 13116 => pixel <= "000000";
      when 13117 => pixel <= "000000";
      when 13118 => pixel <= "000000";
      when 13119 => pixel <= "000000";
      when 13120 => pixel <= "000000";
      when 13121 => pixel <= "000000";
      when 13122 => pixel <= "000000";
      when 13123 => pixel <= "000000";
      when 13124 => pixel <= "000000";
      when 13125 => pixel <= "000000";
      when 13126 => pixel <= "000000";
      when 13127 => pixel <= "000000";
      when 13128 => pixel <= "000000";
      when 13129 => pixel <= "000000";
      when 13130 => pixel <= "000000";
      when 13131 => pixel <= "000000";
      when 13132 => pixel <= "000000";
      when 13133 => pixel <= "000000";
      when 13134 => pixel <= "000000";
      when 13135 => pixel <= "000000";
      when 13136 => pixel <= "000000";
      when 13137 => pixel <= "000000";
      when 13138 => pixel <= "000000";
      when 13139 => pixel <= "000000";
      when 13140 => pixel <= "000000";
      when 13141 => pixel <= "000000";
      when 13142 => pixel <= "000000";
      when 13143 => pixel <= "000000";
      when 13144 => pixel <= "000000";
      when 13145 => pixel <= "000000";
      when 13146 => pixel <= "000000";
      when 13147 => pixel <= "000000";
      when 13148 => pixel <= "000000";
      when 13149 => pixel <= "000000";
      when 13150 => pixel <= "000000";
      when 13151 => pixel <= "000000";
      when 13152 => pixel <= "000000";
      when 13153 => pixel <= "000000";
      when 13154 => pixel <= "000000";
      when 13155 => pixel <= "000000";
      when 13156 => pixel <= "000000";
      when 13157 => pixel <= "000000";
      when 13158 => pixel <= "000000";
      when 13159 => pixel <= "000000";
      when 13160 => pixel <= "000000";
      when 13161 => pixel <= "000000";
      when 13162 => pixel <= "000000";
      when 13163 => pixel <= "000000";
      when 13164 => pixel <= "000000";
      when 13165 => pixel <= "000000";
      when 13166 => pixel <= "000000";
      when 13167 => pixel <= "000000";
      when 13168 => pixel <= "000000";
      when 13169 => pixel <= "000000";
      when 13170 => pixel <= "000000";
      when 13171 => pixel <= "000000";
      when 13172 => pixel <= "000000";
      when 13173 => pixel <= "000000";
      when 13174 => pixel <= "000000";
      when 13175 => pixel <= "000000";
      when 13176 => pixel <= "000000";
      when 13177 => pixel <= "000000";
      when 13178 => pixel <= "000000";
      when 13179 => pixel <= "000000";
      when 13180 => pixel <= "000000";
      when 13181 => pixel <= "000000";
      when 13182 => pixel <= "000000";
      when 13183 => pixel <= "000000";
      when 13184 => pixel <= "000000";
      when 13185 => pixel <= "000000";
      when 13186 => pixel <= "000000";
      when 13187 => pixel <= "000000";
      when 13188 => pixel <= "000000";
      when 13189 => pixel <= "000000";
      when 13190 => pixel <= "000000";
      when 13191 => pixel <= "000000";
      when 13192 => pixel <= "000000";
      when 13193 => pixel <= "000000";
      when 13194 => pixel <= "000000";
      when 13195 => pixel <= "000000";
      when 13196 => pixel <= "000000";
      when 13197 => pixel <= "000000";
      when 13198 => pixel <= "000000";
      when 13199 => pixel <= "000000";
      when 13200 => pixel <= "000000";
      when 13201 => pixel <= "000000";
      when 13202 => pixel <= "000000";
      when 13203 => pixel <= "000000";
      when 13204 => pixel <= "000000";
      when 13205 => pixel <= "000000";
      when 13206 => pixel <= "000000";
      when 13207 => pixel <= "000000";
      when 13208 => pixel <= "000000";
      when 13209 => pixel <= "000000";
      when 13210 => pixel <= "000000";
      when 13211 => pixel <= "000000";
      when 13212 => pixel <= "000000";
      when 13213 => pixel <= "000000";
      when 13214 => pixel <= "000000";
      when 13215 => pixel <= "000000";
      when 13216 => pixel <= "000000";
      when 13217 => pixel <= "000000";
      when 13218 => pixel <= "000000";
      when 13219 => pixel <= "000000";
      when 13220 => pixel <= "000000";
      when 13221 => pixel <= "000000";
      when 13222 => pixel <= "000000";
      when 13223 => pixel <= "000000";
      when 13224 => pixel <= "000000";
      when 13225 => pixel <= "000000";
      when 13226 => pixel <= "000000";
      when 13227 => pixel <= "000000";
      when 13228 => pixel <= "000000";
      when 13229 => pixel <= "000000";
      when 13230 => pixel <= "000000";
      when 13231 => pixel <= "000000";
      when 13232 => pixel <= "000000";
      when 13233 => pixel <= "000000";
      when 13234 => pixel <= "000000";
      when 13235 => pixel <= "000000";
      when 13236 => pixel <= "000000";
      when 13237 => pixel <= "000000";
      when 13238 => pixel <= "000000";
      when 13239 => pixel <= "000000";
      when 13240 => pixel <= "000000";
      when 13241 => pixel <= "000000";
      when 13242 => pixel <= "000000";
      when 13243 => pixel <= "000000";
      when 13244 => pixel <= "000000";
      when 13245 => pixel <= "000000";
      when 13246 => pixel <= "000000";
      when 13247 => pixel <= "000000";
      when 13248 => pixel <= "000000";
      when 13249 => pixel <= "000000";
      when 13250 => pixel <= "000000";
      when 13251 => pixel <= "000000";
      when 13252 => pixel <= "000000";
      when 13253 => pixel <= "000000";
      when 13254 => pixel <= "000000";
      when 13255 => pixel <= "000000";
      when 13256 => pixel <= "000000";
      when 13257 => pixel <= "000000";
      when 13258 => pixel <= "000000";
      when 13259 => pixel <= "000000";
      when 13260 => pixel <= "000000";
      when 13261 => pixel <= "000000";
      when 13262 => pixel <= "000000";
      when 13263 => pixel <= "000000";
      when 13264 => pixel <= "000000";
      when 13265 => pixel <= "000000";
      when 13266 => pixel <= "000000";
      when 13267 => pixel <= "000000";
      when 13268 => pixel <= "000000";
      when 13269 => pixel <= "000000";
      when 13270 => pixel <= "000000";
      when 13271 => pixel <= "000000";
      when 13272 => pixel <= "000000";
      when 13273 => pixel <= "000000";
      when 13274 => pixel <= "000000";
      when 13275 => pixel <= "000000";
      when 13276 => pixel <= "000000";
      when 13277 => pixel <= "000000";
      when 13278 => pixel <= "000000";
      when 13279 => pixel <= "000000";
      when 13280 => pixel <= "000000";
      when 13281 => pixel <= "000000";
      when 13282 => pixel <= "000000";
      when 13283 => pixel <= "000000";
      when 13284 => pixel <= "000000";
      when 13285 => pixel <= "000000";
      when 13286 => pixel <= "000000";
      when 13287 => pixel <= "000000";
      when 13288 => pixel <= "000000";
      when 13289 => pixel <= "000000";
      when 13290 => pixel <= "000000";
      when 13291 => pixel <= "000000";
      when 13292 => pixel <= "000000";
      when 13293 => pixel <= "000000";
      when 13294 => pixel <= "000000";
      when 13295 => pixel <= "000000";
      when 13296 => pixel <= "000000";
      when 13297 => pixel <= "000000";
      when 13298 => pixel <= "000000";
      when 13299 => pixel <= "000000";
      when 13300 => pixel <= "000000";
      when 13301 => pixel <= "000000";
      when 13302 => pixel <= "000000";
      when 13303 => pixel <= "000000";
      when 13304 => pixel <= "000000";
      when 13305 => pixel <= "000000";
      when 13306 => pixel <= "000000";
      when 13307 => pixel <= "000000";
      when 13308 => pixel <= "000000";
      when 13309 => pixel <= "000000";
      when 13310 => pixel <= "000000";
      when 13311 => pixel <= "000000";
      when 13312 => pixel <= "000000";
      when 13313 => pixel <= "000000";
      when 13314 => pixel <= "000000";
      when 13315 => pixel <= "000000";
      when 13316 => pixel <= "000000";
      when 13317 => pixel <= "000000";
      when 13318 => pixel <= "000000";
      when 13319 => pixel <= "000000";
      when 13320 => pixel <= "000000";
      when 13321 => pixel <= "000000";
      when 13322 => pixel <= "000000";
      when 13323 => pixel <= "000000";
      when 13324 => pixel <= "000000";
      when 13325 => pixel <= "000000";
      when 13326 => pixel <= "000000";
      when 13327 => pixel <= "000000";
      when 13328 => pixel <= "000000";
      when 13329 => pixel <= "000000";
      when 13330 => pixel <= "000000";
      when 13331 => pixel <= "000000";
      when 13332 => pixel <= "000000";
      when 13333 => pixel <= "000000";
      when 13334 => pixel <= "000000";
      when 13335 => pixel <= "000000";
      when 13336 => pixel <= "000000";
      when 13337 => pixel <= "000000";
      when 13338 => pixel <= "000000";
      when 13339 => pixel <= "000000";
      when 13340 => pixel <= "000000";
      when 13341 => pixel <= "000000";
      when 13342 => pixel <= "000000";
      when 13343 => pixel <= "000000";
      when 13344 => pixel <= "000000";
      when 13345 => pixel <= "000000";
      when 13346 => pixel <= "000000";
      when 13347 => pixel <= "000000";
      when 13348 => pixel <= "000000";
      when 13349 => pixel <= "000000";
      when 13350 => pixel <= "000000";
      when 13351 => pixel <= "000000";
      when 13352 => pixel <= "000000";
      when 13353 => pixel <= "000000";
      when 13354 => pixel <= "000000";
      when 13355 => pixel <= "000000";
      when 13356 => pixel <= "000000";
      when 13357 => pixel <= "000000";
      when 13358 => pixel <= "000000";
      when 13359 => pixel <= "000000";
      when 13360 => pixel <= "000000";
      when 13361 => pixel <= "000000";
      when 13362 => pixel <= "000000";
      when 13363 => pixel <= "000000";
      when 13364 => pixel <= "000000";
      when 13365 => pixel <= "000000";
      when 13366 => pixel <= "000000";
      when 13367 => pixel <= "000000";
      when 13368 => pixel <= "000000";
      when 13369 => pixel <= "000000";
      when 13370 => pixel <= "000000";
      when 13371 => pixel <= "000000";
      when 13372 => pixel <= "000000";
      when 13373 => pixel <= "000000";
      when 13374 => pixel <= "000000";
      when 13375 => pixel <= "000000";
      when 13376 => pixel <= "000000";
      when 13377 => pixel <= "000000";
      when 13378 => pixel <= "000000";
      when 13379 => pixel <= "000000";
      when 13380 => pixel <= "000000";
      when 13381 => pixel <= "000000";
      when 13382 => pixel <= "000000";
      when 13383 => pixel <= "000000";
      when 13384 => pixel <= "000000";
      when 13385 => pixel <= "000000";
      when 13386 => pixel <= "000000";
      when 13387 => pixel <= "000000";
      when 13388 => pixel <= "000000";
      when 13389 => pixel <= "000000";
      when 13390 => pixel <= "000000";
      when 13391 => pixel <= "000000";
      when 13392 => pixel <= "000000";
      when 13393 => pixel <= "000000";
      when 13394 => pixel <= "000000";
      when 13395 => pixel <= "000000";
      when 13396 => pixel <= "000000";
      when 13397 => pixel <= "000000";
      when 13398 => pixel <= "000000";
      when 13399 => pixel <= "000000";
      when 13400 => pixel <= "000000";
      when 13401 => pixel <= "000000";
      when 13402 => pixel <= "000000";
      when 13403 => pixel <= "000000";
      when 13404 => pixel <= "000000";
      when 13405 => pixel <= "000000";
      when 13406 => pixel <= "000000";
      when 13407 => pixel <= "000000";
      when 13408 => pixel <= "000000";
      when 13409 => pixel <= "000000";
      when 13410 => pixel <= "000000";
      when 13411 => pixel <= "000000";
      when 13412 => pixel <= "000000";
      when 13413 => pixel <= "000000";
      when 13414 => pixel <= "000000";
      when 13415 => pixel <= "000000";
      when 13416 => pixel <= "000000";
      when 13417 => pixel <= "000000";
      when 13418 => pixel <= "000000";
      when 13419 => pixel <= "000000";
      when 13420 => pixel <= "000000";
      when 13421 => pixel <= "000000";
      when 13422 => pixel <= "000000";
      when 13423 => pixel <= "000000";
      when 13424 => pixel <= "000000";
      when 13425 => pixel <= "000000";
      when 13426 => pixel <= "000000";
      when 13427 => pixel <= "000000";
      when 13428 => pixel <= "000000";
      when 13429 => pixel <= "000000";
      when 13430 => pixel <= "000000";
      when 13431 => pixel <= "000000";
      when 13432 => pixel <= "000000";
      when 13433 => pixel <= "000000";
      when 13434 => pixel <= "000000";
      when 13435 => pixel <= "000000";
      when 13436 => pixel <= "000000";
      when 13437 => pixel <= "000000";
      when 13438 => pixel <= "000000";
      when 13439 => pixel <= "000000";
      when 13440 => pixel <= "000000";
      when 13441 => pixel <= "000000";
      when 13442 => pixel <= "000000";
      when 13443 => pixel <= "000000";
      when 13444 => pixel <= "000000";
      when 13445 => pixel <= "000000";
      when 13446 => pixel <= "000000";
      when 13447 => pixel <= "000000";
      when 13448 => pixel <= "000000";
      when 13449 => pixel <= "000000";
      when 13450 => pixel <= "000000";
      when 13451 => pixel <= "000000";
      when 13452 => pixel <= "000000";
      when 13453 => pixel <= "000000";
      when 13454 => pixel <= "000000";
      when 13455 => pixel <= "000000";
      when 13456 => pixel <= "000000";
      when 13457 => pixel <= "000000";
      when 13458 => pixel <= "000000";
      when 13459 => pixel <= "000000";
      when 13460 => pixel <= "000000";
      when 13461 => pixel <= "000000";
      when 13462 => pixel <= "000000";
      when 13463 => pixel <= "000000";
      when 13464 => pixel <= "000000";
      when 13465 => pixel <= "000000";
      when 13466 => pixel <= "000000";
      when 13467 => pixel <= "000000";
      when 13468 => pixel <= "000000";
      when 13469 => pixel <= "000000";
      when 13470 => pixel <= "000000";
      when 13471 => pixel <= "000000";
      when 13472 => pixel <= "000000";
      when 13473 => pixel <= "000000";
      when 13474 => pixel <= "000000";
      when 13475 => pixel <= "000000";
      when 13476 => pixel <= "000000";
      when 13477 => pixel <= "000000";
      when 13478 => pixel <= "000000";
      when 13479 => pixel <= "000000";
      when 13480 => pixel <= "000000";
      when 13481 => pixel <= "000000";
      when 13482 => pixel <= "000000";
      when 13483 => pixel <= "000000";
      when 13484 => pixel <= "000000";
      when 13485 => pixel <= "000000";
      when 13486 => pixel <= "000000";
      when 13487 => pixel <= "000000";
      when 13488 => pixel <= "000000";
      when 13489 => pixel <= "000000";
      when 13490 => pixel <= "000000";
      when 13491 => pixel <= "000000";
      when 13492 => pixel <= "000000";
      when 13493 => pixel <= "000000";
      when 13494 => pixel <= "000000";
      when 13495 => pixel <= "000000";
      when 13496 => pixel <= "000000";
      when 13497 => pixel <= "000000";
      when 13498 => pixel <= "000000";
      when 13499 => pixel <= "000000";
      when 13500 => pixel <= "000000";
      when 13501 => pixel <= "000000";
      when 13502 => pixel <= "000000";
      when 13503 => pixel <= "000000";
      when 13504 => pixel <= "000000";
      when 13505 => pixel <= "000000";
      when 13506 => pixel <= "000000";
      when 13507 => pixel <= "000000";
      when 13508 => pixel <= "000000";
      when 13509 => pixel <= "000000";
      when 13510 => pixel <= "000000";
      when 13511 => pixel <= "000000";
      when 13512 => pixel <= "000000";
      when 13513 => pixel <= "000000";
      when 13514 => pixel <= "000000";
      when 13515 => pixel <= "000000";
      when 13516 => pixel <= "000000";
      when 13517 => pixel <= "000000";
      when 13518 => pixel <= "000000";
      when 13519 => pixel <= "000000";
      when 13520 => pixel <= "000000";
      when 13521 => pixel <= "000000";
      when 13522 => pixel <= "000000";
      when 13523 => pixel <= "000000";
      when 13524 => pixel <= "000000";
      when 13525 => pixel <= "000000";
      when 13526 => pixel <= "000000";
      when 13527 => pixel <= "000000";
      when 13528 => pixel <= "000000";
      when 13529 => pixel <= "000000";
      when 13530 => pixel <= "000000";
      when 13531 => pixel <= "000000";
      when 13532 => pixel <= "000000";
      when 13533 => pixel <= "000000";
      when 13534 => pixel <= "000000";
      when 13535 => pixel <= "000000";
      when 13536 => pixel <= "000000";
      when 13537 => pixel <= "000000";
      when 13538 => pixel <= "000000";
      when 13539 => pixel <= "000000";
      when 13540 => pixel <= "000000";
      when 13541 => pixel <= "000000";
      when 13542 => pixel <= "000000";
      when 13543 => pixel <= "000000";
      when 13544 => pixel <= "000000";
      when 13545 => pixel <= "000000";
      when 13546 => pixel <= "000000";
      when 13547 => pixel <= "000000";
      when 13548 => pixel <= "000000";
      when 13549 => pixel <= "000000";
      when 13550 => pixel <= "000000";
      when 13551 => pixel <= "000000";
      when 13552 => pixel <= "000000";
      when 13553 => pixel <= "000000";
      when 13554 => pixel <= "000000";
      when 13555 => pixel <= "000000";
      when 13556 => pixel <= "000000";
      when 13557 => pixel <= "000000";
      when 13558 => pixel <= "000000";
      when 13559 => pixel <= "000000";
      when 13560 => pixel <= "000000";
      when 13561 => pixel <= "000000";
      when 13562 => pixel <= "000000";
      when 13563 => pixel <= "000000";
      when 13564 => pixel <= "000000";
      when 13565 => pixel <= "000000";
      when 13566 => pixel <= "000000";
      when 13567 => pixel <= "000000";
      when 13568 => pixel <= "000000";
      when 13569 => pixel <= "000000";
      when 13570 => pixel <= "000000";
      when 13571 => pixel <= "000000";
      when 13572 => pixel <= "000000";
      when 13573 => pixel <= "000000";
      when 13574 => pixel <= "000000";
      when 13575 => pixel <= "000000";
      when 13576 => pixel <= "000000";
      when 13577 => pixel <= "000000";
      when 13578 => pixel <= "000000";
      when 13579 => pixel <= "000000";
      when 13580 => pixel <= "000000";
      when 13581 => pixel <= "000000";
      when 13582 => pixel <= "000000";
      when 13583 => pixel <= "000000";
      when 13584 => pixel <= "000000";
      when 13585 => pixel <= "000000";
      when 13586 => pixel <= "000000";
      when 13587 => pixel <= "000000";
      when 13588 => pixel <= "000000";
      when 13589 => pixel <= "000000";
      when 13590 => pixel <= "000000";
      when 13591 => pixel <= "000000";
      when 13592 => pixel <= "000000";
      when 13593 => pixel <= "000000";
      when 13594 => pixel <= "000000";
      when 13595 => pixel <= "000000";
      when 13596 => pixel <= "000000";
      when 13597 => pixel <= "000000";
      when 13598 => pixel <= "000000";
      when 13599 => pixel <= "000000";
      when 13600 => pixel <= "000000";
      when 13601 => pixel <= "000000";
      when 13602 => pixel <= "000000";
      when 13603 => pixel <= "000000";
      when 13604 => pixel <= "000000";
      when 13605 => pixel <= "000000";
      when 13606 => pixel <= "000000";
      when 13607 => pixel <= "000000";
      when 13608 => pixel <= "000000";
      when 13609 => pixel <= "000000";
      when 13610 => pixel <= "000000";
      when 13611 => pixel <= "000000";
      when 13612 => pixel <= "000000";
      when 13613 => pixel <= "000000";
      when 13614 => pixel <= "000000";
      when 13615 => pixel <= "000000";
      when 13616 => pixel <= "000000";
      when 13617 => pixel <= "000000";
      when 13618 => pixel <= "000000";
      when 13619 => pixel <= "000000";
      when 13620 => pixel <= "000000";
      when 13621 => pixel <= "000000";
      when 13622 => pixel <= "000000";
      when 13623 => pixel <= "000000";
      when 13624 => pixel <= "000000";
      when 13625 => pixel <= "000000";
      when 13626 => pixel <= "000000";
      when 13627 => pixel <= "000000";
      when 13628 => pixel <= "000000";
      when 13629 => pixel <= "000000";
      when 13630 => pixel <= "000000";
      when 13631 => pixel <= "000000";
      when 13632 => pixel <= "000000";
      when 13633 => pixel <= "000000";
      when 13634 => pixel <= "000000";
      when 13635 => pixel <= "000000";
      when 13636 => pixel <= "000000";
      when 13637 => pixel <= "000000";
      when 13638 => pixel <= "000000";
      when 13639 => pixel <= "000000";
      when 13640 => pixel <= "000000";
      when 13641 => pixel <= "000000";
      when 13642 => pixel <= "000000";
      when 13643 => pixel <= "000000";
      when 13644 => pixel <= "000000";
      when 13645 => pixel <= "000000";
      when 13646 => pixel <= "000000";
      when 13647 => pixel <= "000000";
      when 13648 => pixel <= "000000";
      when 13649 => pixel <= "000000";
      when 13650 => pixel <= "000000";
      when 13651 => pixel <= "000000";
      when 13652 => pixel <= "000000";
      when 13653 => pixel <= "000000";
      when 13654 => pixel <= "000000";
      when 13655 => pixel <= "000000";
      when 13656 => pixel <= "000000";
      when 13657 => pixel <= "000000";
      when 13658 => pixel <= "000000";
      when 13659 => pixel <= "000000";
      when 13660 => pixel <= "000000";
      when 13661 => pixel <= "000000";
      when 13662 => pixel <= "000000";
      when 13663 => pixel <= "000000";
      when 13664 => pixel <= "000000";
      when 13665 => pixel <= "000000";
      when 13666 => pixel <= "000000";
      when 13667 => pixel <= "000000";
      when 13668 => pixel <= "000000";
      when 13669 => pixel <= "000000";
      when 13670 => pixel <= "000000";
      when 13671 => pixel <= "000000";
      when 13672 => pixel <= "000000";
      when 13673 => pixel <= "000000";
      when 13674 => pixel <= "000000";
      when 13675 => pixel <= "000000";
      when 13676 => pixel <= "000000";
      when 13677 => pixel <= "000000";
      when 13678 => pixel <= "000000";
      when 13679 => pixel <= "000000";
      when 13680 => pixel <= "000000";
      when 13681 => pixel <= "000000";
      when 13682 => pixel <= "000000";
      when 13683 => pixel <= "000000";
      when 13684 => pixel <= "000000";
      when 13685 => pixel <= "000000";
      when 13686 => pixel <= "000000";
      when 13687 => pixel <= "000000";
      when 13688 => pixel <= "000000";
      when 13689 => pixel <= "000000";
      when 13690 => pixel <= "000000";
      when 13691 => pixel <= "000000";
      when 13692 => pixel <= "000000";
      when 13693 => pixel <= "000000";
      when 13694 => pixel <= "000000";
      when 13695 => pixel <= "000000";
      when 13696 => pixel <= "000000";
      when 13697 => pixel <= "000000";
      when 13698 => pixel <= "000000";
      when 13699 => pixel <= "000000";
      when 13700 => pixel <= "000000";
      when 13701 => pixel <= "000000";
      when 13702 => pixel <= "000000";
      when 13703 => pixel <= "000000";
      when 13704 => pixel <= "000000";
      when 13705 => pixel <= "000000";
      when 13706 => pixel <= "000000";
      when 13707 => pixel <= "000000";
      when 13708 => pixel <= "000000";
      when 13709 => pixel <= "000000";
      when 13710 => pixel <= "000000";
      when 13711 => pixel <= "000000";
      when 13712 => pixel <= "000000";
      when 13713 => pixel <= "000000";
      when 13714 => pixel <= "000000";
      when 13715 => pixel <= "000000";
      when 13716 => pixel <= "000000";
      when 13717 => pixel <= "000000";
      when 13718 => pixel <= "000000";
      when 13719 => pixel <= "000000";
      when 13720 => pixel <= "000000";
      when 13721 => pixel <= "000000";
      when 13722 => pixel <= "000000";
      when 13723 => pixel <= "000000";
      when 13724 => pixel <= "000000";
      when 13725 => pixel <= "000000";
      when 13726 => pixel <= "000000";
      when 13727 => pixel <= "000000";
      when 13728 => pixel <= "000000";
      when 13729 => pixel <= "000000";
      when 13730 => pixel <= "000000";
      when 13731 => pixel <= "000000";
      when 13732 => pixel <= "000000";
      when 13733 => pixel <= "000000";
      when 13734 => pixel <= "000000";
      when 13735 => pixel <= "000000";
      when 13736 => pixel <= "000000";
      when 13737 => pixel <= "000000";
      when 13738 => pixel <= "000000";
      when 13739 => pixel <= "000000";
      when 13740 => pixel <= "000000";
      when 13741 => pixel <= "000000";
      when 13742 => pixel <= "000000";
      when 13743 => pixel <= "000000";
      when 13744 => pixel <= "000000";
      when 13745 => pixel <= "000000";
      when 13746 => pixel <= "000000";
      when 13747 => pixel <= "000000";
      when 13748 => pixel <= "000000";
      when 13749 => pixel <= "000000";
      when 13750 => pixel <= "000000";
      when 13751 => pixel <= "000000";
      when 13752 => pixel <= "000000";
      when 13753 => pixel <= "000000";
      when 13754 => pixel <= "000000";
      when 13755 => pixel <= "000000";
      when 13756 => pixel <= "000000";
      when 13757 => pixel <= "000000";
      when 13758 => pixel <= "000000";
      when 13759 => pixel <= "000000";
      when 13760 => pixel <= "000000";
      when 13761 => pixel <= "000000";
      when 13762 => pixel <= "000000";
      when 13763 => pixel <= "000000";
      when 13764 => pixel <= "000000";
      when 13765 => pixel <= "000000";
      when 13766 => pixel <= "000000";
      when 13767 => pixel <= "000000";
      when 13768 => pixel <= "000000";
      when 13769 => pixel <= "000000";
      when 13770 => pixel <= "000000";
      when 13771 => pixel <= "000000";
      when 13772 => pixel <= "000000";
      when 13773 => pixel <= "000000";
      when 13774 => pixel <= "000000";
      when 13775 => pixel <= "000000";
      when 13776 => pixel <= "000000";
      when 13777 => pixel <= "000000";
      when 13778 => pixel <= "000000";
      when 13779 => pixel <= "000000";
      when 13780 => pixel <= "000000";
      when 13781 => pixel <= "000000";
      when 13782 => pixel <= "000000";
      when 13783 => pixel <= "000000";
      when 13784 => pixel <= "000000";
      when 13785 => pixel <= "000000";
      when 13786 => pixel <= "000000";
      when 13787 => pixel <= "000000";
      when 13788 => pixel <= "000000";
      when 13789 => pixel <= "000000";
      when 13790 => pixel <= "000000";
      when 13791 => pixel <= "000000";
      when 13792 => pixel <= "000000";
      when 13793 => pixel <= "000000";
      when 13794 => pixel <= "000000";
      when 13795 => pixel <= "000000";
      when 13796 => pixel <= "000000";
      when 13797 => pixel <= "000000";
      when 13798 => pixel <= "000000";
      when 13799 => pixel <= "000000";
      when 13800 => pixel <= "000000";
      when 13801 => pixel <= "000000";
      when 13802 => pixel <= "000000";
      when 13803 => pixel <= "000000";
      when 13804 => pixel <= "000000";
      when 13805 => pixel <= "000000";
      when 13806 => pixel <= "000000";
      when 13807 => pixel <= "000000";
      when 13808 => pixel <= "000000";
      when 13809 => pixel <= "000000";
      when 13810 => pixel <= "000000";
      when 13811 => pixel <= "000000";
      when 13812 => pixel <= "000000";
      when 13813 => pixel <= "000000";
      when 13814 => pixel <= "000000";
      when 13815 => pixel <= "000000";
      when 13816 => pixel <= "000000";
      when 13817 => pixel <= "000000";
      when 13818 => pixel <= "000000";
      when 13819 => pixel <= "000000";
      when 13820 => pixel <= "000000";
      when 13821 => pixel <= "000000";
      when 13822 => pixel <= "000000";
      when 13823 => pixel <= "000000";
      when 13824 => pixel <= "000000";
      when 13825 => pixel <= "000000";
      when 13826 => pixel <= "000000";
      when 13827 => pixel <= "000000";
      when 13828 => pixel <= "000000";
      when 13829 => pixel <= "000000";
      when 13830 => pixel <= "000000";
      when 13831 => pixel <= "000000";
      when 13832 => pixel <= "000000";
      when 13833 => pixel <= "000000";
      when 13834 => pixel <= "000000";
      when 13835 => pixel <= "000000";
      when 13836 => pixel <= "000000";
      when 13837 => pixel <= "000000";
      when 13838 => pixel <= "000000";
      when 13839 => pixel <= "000000";
      when 13840 => pixel <= "000000";
      when 13841 => pixel <= "000000";
      when 13842 => pixel <= "000000";
      when 13843 => pixel <= "000000";
      when 13844 => pixel <= "000000";
      when 13845 => pixel <= "000000";
      when 13846 => pixel <= "000000";
      when 13847 => pixel <= "000000";
      when 13848 => pixel <= "000000";
      when 13849 => pixel <= "000000";
      when 13850 => pixel <= "000000";
      when 13851 => pixel <= "000000";
      when 13852 => pixel <= "000000";
      when 13853 => pixel <= "000000";
      when 13854 => pixel <= "000000";
      when 13855 => pixel <= "000000";
      when 13856 => pixel <= "000000";
      when 13857 => pixel <= "000000";
      when 13858 => pixel <= "000000";
      when 13859 => pixel <= "000000";
      when 13860 => pixel <= "000000";
      when 13861 => pixel <= "000000";
      when 13862 => pixel <= "000000";
      when 13863 => pixel <= "000000";
      when 13864 => pixel <= "000000";
      when 13865 => pixel <= "000000";
      when 13866 => pixel <= "000000";
      when 13867 => pixel <= "000000";
      when 13868 => pixel <= "000000";
      when 13869 => pixel <= "000000";
      when 13870 => pixel <= "000000";
      when 13871 => pixel <= "000000";
      when 13872 => pixel <= "000000";
      when 13873 => pixel <= "000000";
      when 13874 => pixel <= "000000";
      when 13875 => pixel <= "000000";
      when 13876 => pixel <= "000000";
      when 13877 => pixel <= "000000";
      when 13878 => pixel <= "000000";
      when 13879 => pixel <= "000000";
      when 13880 => pixel <= "000000";
      when 13881 => pixel <= "000000";
      when 13882 => pixel <= "000000";
      when 13883 => pixel <= "000000";
      when 13884 => pixel <= "000000";
      when 13885 => pixel <= "000000";
      when 13886 => pixel <= "000000";
      when 13887 => pixel <= "000000";
      when 13888 => pixel <= "000000";
      when 13889 => pixel <= "000000";
      when 13890 => pixel <= "000000";
      when 13891 => pixel <= "000000";
      when 13892 => pixel <= "000000";
      when 13893 => pixel <= "000000";
      when 13894 => pixel <= "000000";
      when 13895 => pixel <= "000000";
      when 13896 => pixel <= "000000";
      when 13897 => pixel <= "000000";
      when 13898 => pixel <= "000000";
      when 13899 => pixel <= "000000";
      when 13900 => pixel <= "000000";
      when 13901 => pixel <= "000000";
      when 13902 => pixel <= "000000";
      when 13903 => pixel <= "000000";
      when 13904 => pixel <= "000000";
      when 13905 => pixel <= "000000";
      when 13906 => pixel <= "000000";
      when 13907 => pixel <= "000000";
      when 13908 => pixel <= "000000";
      when 13909 => pixel <= "000000";
      when 13910 => pixel <= "000000";
      when 13911 => pixel <= "000000";
      when 13912 => pixel <= "000000";
      when 13913 => pixel <= "000000";
      when 13914 => pixel <= "000000";
      when 13915 => pixel <= "000000";
      when 13916 => pixel <= "000000";
      when 13917 => pixel <= "000000";
      when 13918 => pixel <= "000000";
      when 13919 => pixel <= "000000";
      when 13920 => pixel <= "000000";
      when 13921 => pixel <= "000000";
      when 13922 => pixel <= "000000";
      when 13923 => pixel <= "000000";
      when 13924 => pixel <= "000000";
      when 13925 => pixel <= "000000";
      when 13926 => pixel <= "000000";
      when 13927 => pixel <= "000000";
      when 13928 => pixel <= "000000";
      when 13929 => pixel <= "000000";
      when 13930 => pixel <= "000000";
      when 13931 => pixel <= "000000";
      when 13932 => pixel <= "000000";
      when 13933 => pixel <= "000000";
      when 13934 => pixel <= "000000";
      when 13935 => pixel <= "000000";
      when 13936 => pixel <= "000000";
      when 13937 => pixel <= "000000";
      when 13938 => pixel <= "000000";
      when 13939 => pixel <= "000000";
      when 13940 => pixel <= "000000";
      when 13941 => pixel <= "000000";
      when 13942 => pixel <= "000000";
      when 13943 => pixel <= "000000";
      when 13944 => pixel <= "000000";
      when 13945 => pixel <= "000000";
      when 13946 => pixel <= "000000";
      when 13947 => pixel <= "000000";
      when 13948 => pixel <= "000000";
      when 13949 => pixel <= "000000";
      when 13950 => pixel <= "000000";
      when 13951 => pixel <= "000000";
      when 13952 => pixel <= "000000";
      when 13953 => pixel <= "000000";
      when 13954 => pixel <= "000000";
      when 13955 => pixel <= "000000";
      when 13956 => pixel <= "000000";
      when 13957 => pixel <= "000000";
      when 13958 => pixel <= "000000";
      when 13959 => pixel <= "000000";
      when 13960 => pixel <= "000000";
      when 13961 => pixel <= "000000";
      when 13962 => pixel <= "000000";
      when 13963 => pixel <= "000000";
      when 13964 => pixel <= "000000";
      when 13965 => pixel <= "000000";
      when 13966 => pixel <= "000000";
      when 13967 => pixel <= "000000";
      when 13968 => pixel <= "000000";
      when 13969 => pixel <= "000000";
      when 13970 => pixel <= "000000";
      when 13971 => pixel <= "000000";
      when 13972 => pixel <= "000000";
      when 13973 => pixel <= "000000";
      when 13974 => pixel <= "000000";
      when 13975 => pixel <= "000000";
      when 13976 => pixel <= "000000";
      when 13977 => pixel <= "000000";
      when 13978 => pixel <= "000000";
      when 13979 => pixel <= "000000";
      when 13980 => pixel <= "000000";
      when 13981 => pixel <= "000000";
      when 13982 => pixel <= "000000";
      when 13983 => pixel <= "000000";
      when 13984 => pixel <= "000000";
      when 13985 => pixel <= "000000";
      when 13986 => pixel <= "000000";
      when 13987 => pixel <= "000000";
      when 13988 => pixel <= "000000";
      when 13989 => pixel <= "000000";
      when 13990 => pixel <= "000000";
      when 13991 => pixel <= "000000";
      when 13992 => pixel <= "000000";
      when 13993 => pixel <= "000000";
      when 13994 => pixel <= "000000";
      when 13995 => pixel <= "000000";
      when 13996 => pixel <= "000000";
      when 13997 => pixel <= "000000";
      when 13998 => pixel <= "000000";
      when 13999 => pixel <= "000000";
      when 14000 => pixel <= "000000";
      when 14001 => pixel <= "000000";
      when 14002 => pixel <= "000000";
      when 14003 => pixel <= "000000";
      when 14004 => pixel <= "000000";
      when 14005 => pixel <= "000000";
      when 14006 => pixel <= "000000";
      when 14007 => pixel <= "000000";
      when 14008 => pixel <= "000000";
      when 14009 => pixel <= "000000";
      when 14010 => pixel <= "000000";
      when 14011 => pixel <= "000000";
      when 14012 => pixel <= "000000";
      when 14013 => pixel <= "000000";
      when 14014 => pixel <= "000000";
      when 14015 => pixel <= "000000";
      when 14016 => pixel <= "000000";
      when 14017 => pixel <= "000000";
      when 14018 => pixel <= "000000";
      when 14019 => pixel <= "000000";
      when 14020 => pixel <= "000000";
      when 14021 => pixel <= "000000";
      when 14022 => pixel <= "000000";
      when 14023 => pixel <= "000000";
      when 14024 => pixel <= "000000";
      when 14025 => pixel <= "000000";
      when 14026 => pixel <= "000000";
      when 14027 => pixel <= "000000";
      when 14028 => pixel <= "000000";
      when 14029 => pixel <= "000000";
      when 14030 => pixel <= "000000";
      when 14031 => pixel <= "000000";
      when 14032 => pixel <= "000000";
      when 14033 => pixel <= "000000";
      when 14034 => pixel <= "000000";
      when 14035 => pixel <= "000000";
      when 14036 => pixel <= "000000";
      when 14037 => pixel <= "000000";
      when 14038 => pixel <= "000000";
      when 14039 => pixel <= "000000";
      when 14040 => pixel <= "000000";
      when 14041 => pixel <= "000000";
      when 14042 => pixel <= "000000";
      when 14043 => pixel <= "000000";
      when 14044 => pixel <= "000000";
      when 14045 => pixel <= "000000";
      when 14046 => pixel <= "000000";
      when 14047 => pixel <= "000000";
      when 14048 => pixel <= "000000";
      when 14049 => pixel <= "000000";
      when 14050 => pixel <= "000000";
      when 14051 => pixel <= "000000";
      when 14052 => pixel <= "000000";
      when 14053 => pixel <= "000000";
      when 14054 => pixel <= "000000";
      when 14055 => pixel <= "000000";
      when 14056 => pixel <= "000000";
      when 14057 => pixel <= "000000";
      when 14058 => pixel <= "000000";
      when 14059 => pixel <= "000000";
      when 14060 => pixel <= "000000";
      when 14061 => pixel <= "000000";
      when 14062 => pixel <= "000000";
      when 14063 => pixel <= "000000";
      when 14064 => pixel <= "000000";
      when 14065 => pixel <= "000000";
      when 14066 => pixel <= "000000";
      when 14067 => pixel <= "000000";
      when 14068 => pixel <= "000000";
      when 14069 => pixel <= "000000";
      when 14070 => pixel <= "000000";
      when 14071 => pixel <= "000000";
      when 14072 => pixel <= "000000";
      when 14073 => pixel <= "000000";
      when 14074 => pixel <= "000000";
      when 14075 => pixel <= "000000";
      when 14076 => pixel <= "000000";
      when 14077 => pixel <= "000000";
      when 14078 => pixel <= "000000";
      when 14079 => pixel <= "000000";
      when 14080 => pixel <= "000000";
      when 14081 => pixel <= "000000";
      when 14082 => pixel <= "000000";
      when 14083 => pixel <= "000000";
      when 14084 => pixel <= "000000";
      when 14085 => pixel <= "000000";
      when 14086 => pixel <= "000000";
      when 14087 => pixel <= "000000";
      when 14088 => pixel <= "000000";
      when 14089 => pixel <= "000000";
      when 14090 => pixel <= "000000";
      when 14091 => pixel <= "000000";
      when 14092 => pixel <= "000000";
      when 14093 => pixel <= "000000";
      when 14094 => pixel <= "000000";
      when 14095 => pixel <= "000000";
      when 14096 => pixel <= "000000";
      when 14097 => pixel <= "000000";
      when 14098 => pixel <= "000000";
      when 14099 => pixel <= "000000";
      when 14100 => pixel <= "000000";
      when 14101 => pixel <= "000000";
      when 14102 => pixel <= "000000";
      when 14103 => pixel <= "000000";
      when 14104 => pixel <= "000000";
      when 14105 => pixel <= "000000";
      when 14106 => pixel <= "000000";
      when 14107 => pixel <= "000000";
      when 14108 => pixel <= "000000";
      when 14109 => pixel <= "000000";
      when 14110 => pixel <= "000000";
      when 14111 => pixel <= "000000";
      when 14112 => pixel <= "000000";
      when 14113 => pixel <= "000000";
      when 14114 => pixel <= "000000";
      when 14115 => pixel <= "000000";
      when 14116 => pixel <= "000000";
      when 14117 => pixel <= "000000";
      when 14118 => pixel <= "000000";
      when 14119 => pixel <= "000000";
      when 14120 => pixel <= "000000";
      when 14121 => pixel <= "000000";
      when 14122 => pixel <= "000000";
      when 14123 => pixel <= "000000";
      when 14124 => pixel <= "000000";
      when 14125 => pixel <= "000000";
      when 14126 => pixel <= "000000";
      when 14127 => pixel <= "000000";
      when 14128 => pixel <= "000000";
      when 14129 => pixel <= "000000";
      when 14130 => pixel <= "000000";
      when 14131 => pixel <= "000000";
      when 14132 => pixel <= "000000";
      when 14133 => pixel <= "000000";
      when 14134 => pixel <= "000000";
      when 14135 => pixel <= "000000";
      when 14136 => pixel <= "000000";
      when 14137 => pixel <= "000000";
      when 14138 => pixel <= "000000";
      when 14139 => pixel <= "000000";
      when 14140 => pixel <= "000000";
      when 14141 => pixel <= "000000";
      when 14142 => pixel <= "000000";
      when 14143 => pixel <= "000000";
      when 14144 => pixel <= "000000";
      when 14145 => pixel <= "000000";
      when 14146 => pixel <= "000000";
      when 14147 => pixel <= "000000";
      when 14148 => pixel <= "000000";
      when 14149 => pixel <= "000000";
      when 14150 => pixel <= "000000";
      when 14151 => pixel <= "000000";
      when 14152 => pixel <= "000000";
      when 14153 => pixel <= "000000";
      when 14154 => pixel <= "000000";
      when 14155 => pixel <= "000000";
      when 14156 => pixel <= "000000";
      when 14157 => pixel <= "000000";
      when 14158 => pixel <= "000000";
      when 14159 => pixel <= "000000";
      when 14160 => pixel <= "000000";
      when 14161 => pixel <= "000000";
      when 14162 => pixel <= "000000";
      when 14163 => pixel <= "000000";
      when 14164 => pixel <= "000000";
      when 14165 => pixel <= "000000";
      when 14166 => pixel <= "000000";
      when 14167 => pixel <= "000000";
      when 14168 => pixel <= "000000";
      when 14169 => pixel <= "000000";
      when 14170 => pixel <= "000000";
      when 14171 => pixel <= "000000";
      when 14172 => pixel <= "000000";
      when 14173 => pixel <= "000000";
      when 14174 => pixel <= "000000";
      when 14175 => pixel <= "000000";
      when 14176 => pixel <= "000000";
      when 14177 => pixel <= "000000";
      when 14178 => pixel <= "000000";
      when 14179 => pixel <= "000000";
      when 14180 => pixel <= "000000";
      when 14181 => pixel <= "000000";
      when 14182 => pixel <= "000000";
      when 14183 => pixel <= "000000";
      when 14184 => pixel <= "000000";
      when 14185 => pixel <= "000000";
      when 14186 => pixel <= "000000";
      when 14187 => pixel <= "000000";
      when 14188 => pixel <= "000000";
      when 14189 => pixel <= "000000";
      when 14190 => pixel <= "000000";
      when 14191 => pixel <= "000000";
      when 14192 => pixel <= "000000";
      when 14193 => pixel <= "000000";
      when 14194 => pixel <= "000000";
      when 14195 => pixel <= "000000";
      when 14196 => pixel <= "000000";
      when 14197 => pixel <= "000000";
      when 14198 => pixel <= "000000";
      when 14199 => pixel <= "000000";
      when 14200 => pixel <= "000000";
      when 14201 => pixel <= "000000";
      when 14202 => pixel <= "000000";
      when 14203 => pixel <= "000000";
      when 14204 => pixel <= "000000";
      when 14205 => pixel <= "000000";
      when 14206 => pixel <= "000000";
      when 14207 => pixel <= "000000";
      when 14208 => pixel <= "000000";
      when 14209 => pixel <= "000000";
      when 14210 => pixel <= "000000";
      when 14211 => pixel <= "000000";
      when 14212 => pixel <= "000000";
      when 14213 => pixel <= "000000";
      when 14214 => pixel <= "000000";
      when 14215 => pixel <= "000000";
      when 14216 => pixel <= "000000";
      when 14217 => pixel <= "000000";
      when 14218 => pixel <= "000000";
      when 14219 => pixel <= "000000";
      when 14220 => pixel <= "000000";
      when 14221 => pixel <= "000000";
      when 14222 => pixel <= "000000";
      when 14223 => pixel <= "000000";
      when 14224 => pixel <= "000000";
      when 14225 => pixel <= "000000";
      when 14226 => pixel <= "000000";
      when 14227 => pixel <= "000000";
      when 14228 => pixel <= "000000";
      when 14229 => pixel <= "000000";
      when 14230 => pixel <= "000000";
      when 14231 => pixel <= "000000";
      when 14232 => pixel <= "000000";
      when 14233 => pixel <= "000000";
      when 14234 => pixel <= "000000";
      when 14235 => pixel <= "000000";
      when 14236 => pixel <= "000000";
      when 14237 => pixel <= "000000";
      when 14238 => pixel <= "000000";
      when 14239 => pixel <= "000000";
      when 14240 => pixel <= "000000";
      when 14241 => pixel <= "000000";
      when 14242 => pixel <= "000000";
      when 14243 => pixel <= "000000";
      when 14244 => pixel <= "000000";
      when 14245 => pixel <= "000000";
      when 14246 => pixel <= "000000";
      when 14247 => pixel <= "000000";
      when 14248 => pixel <= "000000";
      when 14249 => pixel <= "000000";
      when 14250 => pixel <= "000000";
      when 14251 => pixel <= "000000";
      when 14252 => pixel <= "000000";
      when 14253 => pixel <= "000000";
      when 14254 => pixel <= "000000";
      when 14255 => pixel <= "000000";
      when 14256 => pixel <= "000000";
      when 14257 => pixel <= "000000";
      when 14258 => pixel <= "000000";
      when 14259 => pixel <= "000000";
      when 14260 => pixel <= "000000";
      when 14261 => pixel <= "000000";
      when 14262 => pixel <= "000000";
      when 14263 => pixel <= "000000";
      when 14264 => pixel <= "000000";
      when 14265 => pixel <= "000000";
      when 14266 => pixel <= "000000";
      when 14267 => pixel <= "000000";
      when 14268 => pixel <= "000000";
      when 14269 => pixel <= "000000";
      when 14270 => pixel <= "000000";
      when 14271 => pixel <= "000000";
      when 14272 => pixel <= "000000";
      when 14273 => pixel <= "000000";
      when 14274 => pixel <= "000000";
      when 14275 => pixel <= "000000";
      when 14276 => pixel <= "000000";
      when 14277 => pixel <= "000000";
      when 14278 => pixel <= "000000";
      when 14279 => pixel <= "000000";
      when 14280 => pixel <= "000000";
      when 14281 => pixel <= "000000";
      when 14282 => pixel <= "000000";
      when 14283 => pixel <= "000000";
      when 14284 => pixel <= "000000";
      when 14285 => pixel <= "000000";
      when 14286 => pixel <= "000000";
      when 14287 => pixel <= "000000";
      when 14288 => pixel <= "000000";
      when 14289 => pixel <= "000000";
      when 14290 => pixel <= "000000";
      when 14291 => pixel <= "000000";
      when 14292 => pixel <= "000000";
      when 14293 => pixel <= "000000";
      when 14294 => pixel <= "000000";
      when 14295 => pixel <= "000000";
      when 14296 => pixel <= "000000";
      when 14297 => pixel <= "000000";
      when 14298 => pixel <= "000000";
      when 14299 => pixel <= "000000";
      when 14300 => pixel <= "000000";
      when 14301 => pixel <= "000000";
      when 14302 => pixel <= "000000";
      when 14303 => pixel <= "000000";
      when 14304 => pixel <= "000000";
      when 14305 => pixel <= "000000";
      when 14306 => pixel <= "000000";
      when 14307 => pixel <= "000000";
      when 14308 => pixel <= "000000";
      when 14309 => pixel <= "000000";
      when 14310 => pixel <= "000000";
      when 14311 => pixel <= "000000";
      when 14312 => pixel <= "000000";
      when 14313 => pixel <= "000000";
      when 14314 => pixel <= "000000";
      when 14315 => pixel <= "000000";
      when 14316 => pixel <= "000000";
      when 14317 => pixel <= "000000";
      when 14318 => pixel <= "000000";
      when 14319 => pixel <= "000000";
      when 14320 => pixel <= "000000";
      when 14321 => pixel <= "000000";
      when 14322 => pixel <= "000000";
      when 14323 => pixel <= "000000";
      when 14324 => pixel <= "000000";
      when 14325 => pixel <= "000000";
      when 14326 => pixel <= "000000";
      when 14327 => pixel <= "000000";
      when 14328 => pixel <= "000000";
      when 14329 => pixel <= "000000";
      when 14330 => pixel <= "000000";
      when 14331 => pixel <= "000000";
      when 14332 => pixel <= "000000";
      when 14333 => pixel <= "000000";
      when 14334 => pixel <= "000000";
      when 14335 => pixel <= "000000";
      when 14336 => pixel <= "000000";
      when 14337 => pixel <= "000000";
      when 14338 => pixel <= "000000";
      when 14339 => pixel <= "000000";
      when 14340 => pixel <= "000000";
      when 14341 => pixel <= "000000";
      when 14342 => pixel <= "000000";
      when 14343 => pixel <= "000000";
      when 14344 => pixel <= "000000";
      when 14345 => pixel <= "000000";
      when 14346 => pixel <= "000000";
      when 14347 => pixel <= "000000";
      when 14348 => pixel <= "000000";
      when 14349 => pixel <= "000000";
      when 14350 => pixel <= "000000";
      when 14351 => pixel <= "000000";
      when 14352 => pixel <= "000000";
      when 14353 => pixel <= "000000";
      when 14354 => pixel <= "000000";
      when 14355 => pixel <= "000000";
      when 14356 => pixel <= "000000";
      when 14357 => pixel <= "000000";
      when 14358 => pixel <= "000000";
      when 14359 => pixel <= "000000";
      when 14360 => pixel <= "000000";
      when 14361 => pixel <= "000000";
      when 14362 => pixel <= "000000";
      when 14363 => pixel <= "000000";
      when 14364 => pixel <= "000000";
      when 14365 => pixel <= "000000";
      when 14366 => pixel <= "000000";
      when 14367 => pixel <= "000000";
      when 14368 => pixel <= "000000";
      when 14369 => pixel <= "000000";
      when 14370 => pixel <= "000000";
      when 14371 => pixel <= "000000";
      when 14372 => pixel <= "000000";
      when 14373 => pixel <= "000000";
      when 14374 => pixel <= "000000";
      when 14375 => pixel <= "000000";
      when 14376 => pixel <= "000000";
      when 14377 => pixel <= "000000";
      when 14378 => pixel <= "000000";
      when 14379 => pixel <= "000000";
      when 14380 => pixel <= "000000";
      when 14381 => pixel <= "000000";
      when 14382 => pixel <= "000000";
      when 14383 => pixel <= "000000";
      when 14384 => pixel <= "000000";
      when 14385 => pixel <= "000000";
      when 14386 => pixel <= "000000";
      when 14387 => pixel <= "000000";
      when 14388 => pixel <= "000000";
      when 14389 => pixel <= "000000";
      when 14390 => pixel <= "000000";
      when 14391 => pixel <= "000000";
      when 14392 => pixel <= "000000";
      when 14393 => pixel <= "000000";
      when 14394 => pixel <= "000000";
      when 14395 => pixel <= "000000";
      when 14396 => pixel <= "000000";
      when 14397 => pixel <= "000000";
      when 14398 => pixel <= "000000";
      when 14399 => pixel <= "000000";
      when 14400 => pixel <= "000000";
      when 14401 => pixel <= "000000";
      when 14402 => pixel <= "000000";
      when 14403 => pixel <= "000000";
      when 14404 => pixel <= "000000";
      when 14405 => pixel <= "000000";
      when 14406 => pixel <= "000000";
      when 14407 => pixel <= "000000";
      when 14408 => pixel <= "000000";
      when 14409 => pixel <= "000000";
      when 14410 => pixel <= "000000";
      when 14411 => pixel <= "000000";
      when 14412 => pixel <= "000000";
      when 14413 => pixel <= "000000";
      when 14414 => pixel <= "000000";
      when 14415 => pixel <= "000000";
      when 14416 => pixel <= "000000";
      when 14417 => pixel <= "000000";
      when 14418 => pixel <= "000000";
      when 14419 => pixel <= "000000";
      when 14420 => pixel <= "000000";
      when 14421 => pixel <= "000000";
      when 14422 => pixel <= "000000";
      when 14423 => pixel <= "000000";
      when 14424 => pixel <= "000000";
      when 14425 => pixel <= "000000";
      when 14426 => pixel <= "000000";
      when 14427 => pixel <= "000000";
      when 14428 => pixel <= "000000";
      when 14429 => pixel <= "000000";
      when 14430 => pixel <= "000000";
      when 14431 => pixel <= "000000";
      when 14432 => pixel <= "000000";
      when 14433 => pixel <= "000000";
      when 14434 => pixel <= "000000";
      when 14435 => pixel <= "000000";
      when 14436 => pixel <= "000000";
      when 14437 => pixel <= "000000";
      when 14438 => pixel <= "000000";
      when 14439 => pixel <= "000000";
      when 14440 => pixel <= "000000";
      when 14441 => pixel <= "000000";
      when 14442 => pixel <= "000000";
      when 14443 => pixel <= "000000";
      when 14444 => pixel <= "000000";
      when 14445 => pixel <= "000000";
      when 14446 => pixel <= "000000";
      when 14447 => pixel <= "000000";
      when 14448 => pixel <= "000000";
      when 14449 => pixel <= "000000";
      when 14450 => pixel <= "000000";
      when 14451 => pixel <= "000000";
      when 14452 => pixel <= "000000";
      when 14453 => pixel <= "000000";
      when 14454 => pixel <= "000000";
      when 14455 => pixel <= "000000";
      when 14456 => pixel <= "000000";
      when 14457 => pixel <= "000000";
      when 14458 => pixel <= "000000";
      when 14459 => pixel <= "000000";
      when 14460 => pixel <= "000000";
      when 14461 => pixel <= "000000";
      when 14462 => pixel <= "000000";
      when 14463 => pixel <= "000000";
      when 14464 => pixel <= "000000";
      when 14465 => pixel <= "000000";
      when 14466 => pixel <= "000000";
      when 14467 => pixel <= "000000";
      when 14468 => pixel <= "000000";
      when 14469 => pixel <= "000000";
      when 14470 => pixel <= "000000";
      when 14471 => pixel <= "000000";
      when 14472 => pixel <= "000000";
      when 14473 => pixel <= "000000";
      when 14474 => pixel <= "000000";
      when 14475 => pixel <= "000000";
      when 14476 => pixel <= "000000";
      when 14477 => pixel <= "000000";
      when 14478 => pixel <= "000000";
      when 14479 => pixel <= "000000";
      when 14480 => pixel <= "000000";
      when 14481 => pixel <= "000000";
      when 14482 => pixel <= "000000";
      when 14483 => pixel <= "000000";
      when 14484 => pixel <= "000000";
      when 14485 => pixel <= "000000";
      when 14486 => pixel <= "000000";
      when 14487 => pixel <= "000000";
      when 14488 => pixel <= "000000";
      when 14489 => pixel <= "000000";
      when 14490 => pixel <= "000000";
      when 14491 => pixel <= "000000";
      when 14492 => pixel <= "000000";
      when 14493 => pixel <= "000000";
      when 14494 => pixel <= "000000";
      when 14495 => pixel <= "000000";
      when 14496 => pixel <= "000000";
      when 14497 => pixel <= "000000";
      when 14498 => pixel <= "000000";
      when 14499 => pixel <= "000000";
      when 14500 => pixel <= "000000";
      when 14501 => pixel <= "000000";
      when 14502 => pixel <= "000000";
      when 14503 => pixel <= "000000";
      when 14504 => pixel <= "000000";
      when 14505 => pixel <= "000000";
      when 14506 => pixel <= "000000";
      when 14507 => pixel <= "000000";
      when 14508 => pixel <= "000000";
      when 14509 => pixel <= "000000";
      when 14510 => pixel <= "000000";
      when 14511 => pixel <= "000000";
      when 14512 => pixel <= "000000";
      when 14513 => pixel <= "000000";
      when 14514 => pixel <= "000000";
      when 14515 => pixel <= "000000";
      when 14516 => pixel <= "000000";
      when 14517 => pixel <= "000000";
      when 14518 => pixel <= "000000";
      when 14519 => pixel <= "000000";
      when 14520 => pixel <= "000000";
      when 14521 => pixel <= "000000";
      when 14522 => pixel <= "000000";
      when 14523 => pixel <= "000000";
      when 14524 => pixel <= "000000";
      when 14525 => pixel <= "000000";
      when 14526 => pixel <= "000000";
      when 14527 => pixel <= "000000";
      when 14528 => pixel <= "000000";
      when 14529 => pixel <= "000000";
      when 14530 => pixel <= "000000";
      when 14531 => pixel <= "000000";
      when 14532 => pixel <= "000000";
      when 14533 => pixel <= "000000";
      when 14534 => pixel <= "000000";
      when 14535 => pixel <= "000000";
      when 14536 => pixel <= "000000";
      when 14537 => pixel <= "000000";
      when 14538 => pixel <= "000000";
      when 14539 => pixel <= "000000";
      when 14540 => pixel <= "000000";
      when 14541 => pixel <= "000000";
      when 14542 => pixel <= "000000";
      when 14543 => pixel <= "000000";
      when 14544 => pixel <= "000000";
      when 14545 => pixel <= "000000";
      when 14546 => pixel <= "000000";
      when 14547 => pixel <= "000000";
      when 14548 => pixel <= "000000";
      when 14549 => pixel <= "000000";
      when 14550 => pixel <= "000000";
      when 14551 => pixel <= "000000";
      when 14552 => pixel <= "000000";
      when 14553 => pixel <= "000000";
      when 14554 => pixel <= "000000";
      when 14555 => pixel <= "000000";
      when 14556 => pixel <= "000000";
      when 14557 => pixel <= "000000";
      when 14558 => pixel <= "000000";
      when 14559 => pixel <= "000000";
      when 14560 => pixel <= "000000";
      when 14561 => pixel <= "000000";
      when 14562 => pixel <= "000000";
      when 14563 => pixel <= "000000";
      when 14564 => pixel <= "000000";
      when 14565 => pixel <= "000000";
      when 14566 => pixel <= "000000";
      when 14567 => pixel <= "000000";
      when 14568 => pixel <= "000000";
      when 14569 => pixel <= "000000";
      when 14570 => pixel <= "000000";
      when 14571 => pixel <= "000000";
      when 14572 => pixel <= "000000";
      when 14573 => pixel <= "000000";
      when 14574 => pixel <= "000000";
      when 14575 => pixel <= "000000";
      when 14576 => pixel <= "000000";
      when 14577 => pixel <= "000000";
      when 14578 => pixel <= "000000";
      when 14579 => pixel <= "000000";
      when 14580 => pixel <= "000000";
      when 14581 => pixel <= "000000";
      when 14582 => pixel <= "000000";
      when 14583 => pixel <= "000000";
      when 14584 => pixel <= "000000";
      when 14585 => pixel <= "000000";
      when 14586 => pixel <= "000000";
      when 14587 => pixel <= "000000";
      when 14588 => pixel <= "000000";
      when 14589 => pixel <= "000000";
      when 14590 => pixel <= "000000";
      when 14591 => pixel <= "000000";
      when 14592 => pixel <= "000000";
      when 14593 => pixel <= "000000";
      when 14594 => pixel <= "000000";
      when 14595 => pixel <= "000000";
      when 14596 => pixel <= "000000";
      when 14597 => pixel <= "000000";
      when 14598 => pixel <= "000000";
      when 14599 => pixel <= "000000";
      when 14600 => pixel <= "000000";
      when 14601 => pixel <= "000000";
      when 14602 => pixel <= "000000";
      when 14603 => pixel <= "000000";
      when 14604 => pixel <= "000000";
      when 14605 => pixel <= "000000";
      when 14606 => pixel <= "000000";
      when 14607 => pixel <= "000000";
      when 14608 => pixel <= "000000";
      when 14609 => pixel <= "000000";
      when 14610 => pixel <= "000000";
      when 14611 => pixel <= "000000";
      when 14612 => pixel <= "000000";
      when 14613 => pixel <= "000000";
      when 14614 => pixel <= "000000";
      when 14615 => pixel <= "000000";
      when 14616 => pixel <= "000000";
      when 14617 => pixel <= "000000";
      when 14618 => pixel <= "000000";
      when 14619 => pixel <= "000000";
      when 14620 => pixel <= "000000";
      when 14621 => pixel <= "000000";
      when 14622 => pixel <= "000000";
      when 14623 => pixel <= "000000";
      when 14624 => pixel <= "000000";
      when 14625 => pixel <= "000000";
      when 14626 => pixel <= "000000";
      when 14627 => pixel <= "000000";
      when 14628 => pixel <= "000000";
      when 14629 => pixel <= "000000";
      when 14630 => pixel <= "000000";
      when 14631 => pixel <= "000000";
      when 14632 => pixel <= "000000";
      when 14633 => pixel <= "000000";
      when 14634 => pixel <= "000000";
      when 14635 => pixel <= "000000";
      when 14636 => pixel <= "000000";
      when 14637 => pixel <= "000000";
      when 14638 => pixel <= "000000";
      when 14639 => pixel <= "000000";
      when 14640 => pixel <= "000000";
      when 14641 => pixel <= "000000";
      when 14642 => pixel <= "000000";
      when 14643 => pixel <= "000000";
      when 14644 => pixel <= "000000";
      when 14645 => pixel <= "000000";
      when 14646 => pixel <= "000000";
      when 14647 => pixel <= "000000";
      when 14648 => pixel <= "000000";
      when 14649 => pixel <= "000000";
      when 14650 => pixel <= "000000";
      when 14651 => pixel <= "000000";
      when 14652 => pixel <= "000000";
      when 14653 => pixel <= "000000";
      when 14654 => pixel <= "000000";
      when 14655 => pixel <= "000000";
      when 14656 => pixel <= "000000";
      when 14657 => pixel <= "000000";
      when 14658 => pixel <= "000000";
      when 14659 => pixel <= "000000";
      when 14660 => pixel <= "000000";
      when 14661 => pixel <= "000000";
      when 14662 => pixel <= "000000";
      when 14663 => pixel <= "000000";
      when 14664 => pixel <= "000000";
      when 14665 => pixel <= "000000";
      when 14666 => pixel <= "000000";
      when 14667 => pixel <= "000000";
      when 14668 => pixel <= "000000";
      when 14669 => pixel <= "000000";
      when 14670 => pixel <= "000000";
      when 14671 => pixel <= "000000";
      when 14672 => pixel <= "000000";
      when 14673 => pixel <= "000000";
      when 14674 => pixel <= "000000";
      when 14675 => pixel <= "000000";
      when 14676 => pixel <= "000000";
      when 14677 => pixel <= "000000";
      when 14678 => pixel <= "000000";
      when 14679 => pixel <= "000000";
      when 14680 => pixel <= "000000";
      when 14681 => pixel <= "000000";
      when 14682 => pixel <= "000000";
      when 14683 => pixel <= "000000";
      when 14684 => pixel <= "000000";
      when 14685 => pixel <= "000000";
      when 14686 => pixel <= "000000";
      when 14687 => pixel <= "000000";
      when 14688 => pixel <= "000000";
      when 14689 => pixel <= "000000";
      when 14690 => pixel <= "000000";
      when 14691 => pixel <= "000000";
      when 14692 => pixel <= "000000";
      when 14693 => pixel <= "000000";
      when 14694 => pixel <= "000000";
      when 14695 => pixel <= "000000";
      when 14696 => pixel <= "000000";
      when 14697 => pixel <= "000000";
      when 14698 => pixel <= "000000";
      when 14699 => pixel <= "000000";
      when 14700 => pixel <= "000000";
      when 14701 => pixel <= "000000";
      when 14702 => pixel <= "000000";
      when 14703 => pixel <= "000000";
      when 14704 => pixel <= "000000";
      when 14705 => pixel <= "000000";
      when 14706 => pixel <= "000000";
      when 14707 => pixel <= "000000";
      when 14708 => pixel <= "000000";
      when 14709 => pixel <= "000000";
      when 14710 => pixel <= "000000";
      when 14711 => pixel <= "000000";
      when 14712 => pixel <= "000000";
      when 14713 => pixel <= "000000";
      when 14714 => pixel <= "000000";
      when 14715 => pixel <= "000000";
      when 14716 => pixel <= "000000";
      when 14717 => pixel <= "000000";
      when 14718 => pixel <= "000000";
      when 14719 => pixel <= "000000";
      when 14720 => pixel <= "000000";
      when 14721 => pixel <= "000000";
      when 14722 => pixel <= "000000";
      when 14723 => pixel <= "000000";
      when 14724 => pixel <= "000000";
      when 14725 => pixel <= "000000";
      when 14726 => pixel <= "000000";
      when 14727 => pixel <= "000000";
      when 14728 => pixel <= "000000";
      when 14729 => pixel <= "000000";
      when 14730 => pixel <= "000000";
      when 14731 => pixel <= "000000";
      when 14732 => pixel <= "000000";
      when 14733 => pixel <= "000000";
      when 14734 => pixel <= "000000";
      when 14735 => pixel <= "000000";
      when 14736 => pixel <= "000000";
      when 14737 => pixel <= "000000";
      when 14738 => pixel <= "000000";
      when 14739 => pixel <= "000000";
      when 14740 => pixel <= "000000";
      when 14741 => pixel <= "000000";
      when 14742 => pixel <= "000000";
      when 14743 => pixel <= "000000";
      when 14744 => pixel <= "000000";
      when 14745 => pixel <= "000000";
      when 14746 => pixel <= "000000";
      when 14747 => pixel <= "000000";
      when 14748 => pixel <= "000000";
      when 14749 => pixel <= "000000";
      when 14750 => pixel <= "000000";
      when 14751 => pixel <= "000000";
      when 14752 => pixel <= "000000";
      when 14753 => pixel <= "000000";
      when 14754 => pixel <= "000000";
      when 14755 => pixel <= "000000";
      when 14756 => pixel <= "000000";
      when 14757 => pixel <= "000000";
      when 14758 => pixel <= "000000";
      when 14759 => pixel <= "000000";
      when 14760 => pixel <= "000000";
      when 14761 => pixel <= "000000";
      when 14762 => pixel <= "000000";
      when 14763 => pixel <= "000000";
      when 14764 => pixel <= "000000";
      when 14765 => pixel <= "000000";
      when 14766 => pixel <= "000000";
      when 14767 => pixel <= "000000";
      when 14768 => pixel <= "000000";
      when 14769 => pixel <= "000000";
      when 14770 => pixel <= "000000";
      when 14771 => pixel <= "000000";
      when 14772 => pixel <= "000000";
      when 14773 => pixel <= "000000";
      when 14774 => pixel <= "000000";
      when 14775 => pixel <= "000000";
      when 14776 => pixel <= "000000";
      when 14777 => pixel <= "000000";
      when 14778 => pixel <= "000000";
      when 14779 => pixel <= "000000";
      when 14780 => pixel <= "000000";
      when 14781 => pixel <= "000000";
      when 14782 => pixel <= "000000";
      when 14783 => pixel <= "000000";
      when 14784 => pixel <= "000000";
      when 14785 => pixel <= "000000";
      when 14786 => pixel <= "000000";
      when 14787 => pixel <= "000000";
      when 14788 => pixel <= "000000";
      when 14789 => pixel <= "000000";
      when 14790 => pixel <= "000000";
      when 14791 => pixel <= "000000";
      when 14792 => pixel <= "000000";
      when 14793 => pixel <= "000000";
      when 14794 => pixel <= "000000";
      when 14795 => pixel <= "000000";
      when 14796 => pixel <= "000000";
      when 14797 => pixel <= "000000";
      when 14798 => pixel <= "000000";
      when 14799 => pixel <= "000000";
      when 14800 => pixel <= "000000";
      when 14801 => pixel <= "000000";
      when 14802 => pixel <= "000000";
      when 14803 => pixel <= "000000";
      when 14804 => pixel <= "000000";
      when 14805 => pixel <= "000000";
      when 14806 => pixel <= "000000";
      when 14807 => pixel <= "000000";
      when 14808 => pixel <= "000000";
      when 14809 => pixel <= "000000";
      when 14810 => pixel <= "000000";
      when 14811 => pixel <= "000000";
      when 14812 => pixel <= "000000";
      when 14813 => pixel <= "000000";
      when 14814 => pixel <= "000000";
      when 14815 => pixel <= "000000";
      when 14816 => pixel <= "000000";
      when 14817 => pixel <= "000000";
      when 14818 => pixel <= "000000";
      when 14819 => pixel <= "000000";
      when 14820 => pixel <= "000000";
      when 14821 => pixel <= "000000";
      when 14822 => pixel <= "000000";
      when 14823 => pixel <= "000000";
      when 14824 => pixel <= "000000";
      when 14825 => pixel <= "000000";
      when 14826 => pixel <= "000000";
      when 14827 => pixel <= "000000";
      when 14828 => pixel <= "000000";
      when 14829 => pixel <= "000000";
      when 14830 => pixel <= "000000";
      when 14831 => pixel <= "000000";
      when 14832 => pixel <= "000000";
      when 14833 => pixel <= "000000";
      when 14834 => pixel <= "000000";
      when 14835 => pixel <= "000000";
      when 14836 => pixel <= "000000";
      when 14837 => pixel <= "000000";
      when 14838 => pixel <= "000000";
      when 14839 => pixel <= "000000";
      when 14840 => pixel <= "000000";
      when 14841 => pixel <= "000000";
      when 14842 => pixel <= "000000";
      when 14843 => pixel <= "000000";
      when 14844 => pixel <= "000000";
      when 14845 => pixel <= "000000";
      when 14846 => pixel <= "000000";
      when 14847 => pixel <= "000000";
      when 14848 => pixel <= "000000";
      when 14849 => pixel <= "000000";
      when 14850 => pixel <= "000000";
      when 14851 => pixel <= "000000";
      when 14852 => pixel <= "000000";
      when 14853 => pixel <= "000000";
      when 14854 => pixel <= "000000";
      when 14855 => pixel <= "000000";
      when 14856 => pixel <= "000000";
      when 14857 => pixel <= "000000";
      when 14858 => pixel <= "000000";
      when 14859 => pixel <= "000000";
      when 14860 => pixel <= "000000";
      when 14861 => pixel <= "000000";
      when 14862 => pixel <= "000000";
      when 14863 => pixel <= "000000";
      when 14864 => pixel <= "000000";
      when 14865 => pixel <= "000000";
      when 14866 => pixel <= "000000";
      when 14867 => pixel <= "000000";
      when 14868 => pixel <= "000000";
      when 14869 => pixel <= "000000";
      when 14870 => pixel <= "000000";
      when 14871 => pixel <= "000000";
      when 14872 => pixel <= "000000";
      when 14873 => pixel <= "000000";
      when 14874 => pixel <= "000000";
      when 14875 => pixel <= "000000";
      when 14876 => pixel <= "000000";
      when 14877 => pixel <= "000000";
      when 14878 => pixel <= "000000";
      when 14879 => pixel <= "000000";
      when 14880 => pixel <= "000000";
      when 14881 => pixel <= "000000";
      when 14882 => pixel <= "000000";
      when 14883 => pixel <= "000000";
      when 14884 => pixel <= "000000";
      when 14885 => pixel <= "000000";
      when 14886 => pixel <= "000000";
      when 14887 => pixel <= "000000";
      when 14888 => pixel <= "000000";
      when 14889 => pixel <= "000000";
      when 14890 => pixel <= "000000";
      when 14891 => pixel <= "000000";
      when 14892 => pixel <= "000000";
      when 14893 => pixel <= "000000";
      when 14894 => pixel <= "000000";
      when 14895 => pixel <= "000000";
      when 14896 => pixel <= "000000";
      when 14897 => pixel <= "000000";
      when 14898 => pixel <= "000000";
      when 14899 => pixel <= "000000";
      when 14900 => pixel <= "000000";
      when 14901 => pixel <= "000000";
      when 14902 => pixel <= "000000";
      when 14903 => pixel <= "000000";
      when 14904 => pixel <= "000000";
      when 14905 => pixel <= "000000";
      when 14906 => pixel <= "000000";
      when 14907 => pixel <= "000000";
      when 14908 => pixel <= "000000";
      when 14909 => pixel <= "000000";
      when 14910 => pixel <= "000000";
      when 14911 => pixel <= "000000";
      when 14912 => pixel <= "000000";
      when 14913 => pixel <= "000000";
      when 14914 => pixel <= "000000";
      when 14915 => pixel <= "000000";
      when 14916 => pixel <= "000000";
      when 14917 => pixel <= "000000";
      when 14918 => pixel <= "000000";
      when 14919 => pixel <= "000000";
      when 14920 => pixel <= "000000";
      when 14921 => pixel <= "000000";
      when 14922 => pixel <= "000000";
      when 14923 => pixel <= "000000";
      when 14924 => pixel <= "000000";
      when 14925 => pixel <= "000000";
      when 14926 => pixel <= "000000";
      when 14927 => pixel <= "000000";
      when 14928 => pixel <= "000000";
      when 14929 => pixel <= "000000";
      when 14930 => pixel <= "000000";
      when 14931 => pixel <= "000000";
      when 14932 => pixel <= "000000";
      when 14933 => pixel <= "000000";
      when 14934 => pixel <= "000000";
      when 14935 => pixel <= "000000";
      when 14936 => pixel <= "000000";
      when 14937 => pixel <= "000000";
      when 14938 => pixel <= "000000";
      when 14939 => pixel <= "000000";
      when 14940 => pixel <= "000000";
      when 14941 => pixel <= "000000";
      when 14942 => pixel <= "000000";
      when 14943 => pixel <= "000000";
      when 14944 => pixel <= "000000";
      when 14945 => pixel <= "000000";
      when 14946 => pixel <= "000000";
      when 14947 => pixel <= "000000";
      when 14948 => pixel <= "000000";
      when 14949 => pixel <= "000000";
      when 14950 => pixel <= "000000";
      when 14951 => pixel <= "000000";
      when 14952 => pixel <= "000000";
      when 14953 => pixel <= "000000";
      when 14954 => pixel <= "000000";
      when 14955 => pixel <= "000000";
      when 14956 => pixel <= "000000";
      when 14957 => pixel <= "000000";
      when 14958 => pixel <= "000000";
      when 14959 => pixel <= "000000";
      when 14960 => pixel <= "000000";
      when 14961 => pixel <= "000000";
      when 14962 => pixel <= "000000";
      when 14963 => pixel <= "000000";
      when 14964 => pixel <= "000000";
      when 14965 => pixel <= "000000";
      when 14966 => pixel <= "000000";
      when 14967 => pixel <= "000000";
      when 14968 => pixel <= "000000";
      when 14969 => pixel <= "000000";
      when 14970 => pixel <= "000000";
      when 14971 => pixel <= "000000";
      when 14972 => pixel <= "000000";
      when 14973 => pixel <= "000000";
      when 14974 => pixel <= "000000";
      when 14975 => pixel <= "000000";
      when 14976 => pixel <= "000000";
      when 14977 => pixel <= "000000";
      when 14978 => pixel <= "000000";
      when 14979 => pixel <= "000000";
      when 14980 => pixel <= "000000";
      when 14981 => pixel <= "000000";
      when 14982 => pixel <= "000000";
      when 14983 => pixel <= "000000";
      when 14984 => pixel <= "000000";
      when 14985 => pixel <= "000000";
      when 14986 => pixel <= "000000";
      when 14987 => pixel <= "000000";
      when 14988 => pixel <= "000000";
      when 14989 => pixel <= "000000";
      when 14990 => pixel <= "000000";
      when 14991 => pixel <= "000000";
      when 14992 => pixel <= "000000";
      when 14993 => pixel <= "000000";
      when 14994 => pixel <= "000000";
      when 14995 => pixel <= "000000";
      when 14996 => pixel <= "000000";
      when 14997 => pixel <= "000000";
      when 14998 => pixel <= "000000";
      when 14999 => pixel <= "000000";
      when 15000 => pixel <= "000000";
      when 15001 => pixel <= "000000";
      when 15002 => pixel <= "000000";
      when 15003 => pixel <= "000000";
      when 15004 => pixel <= "000000";
      when 15005 => pixel <= "000000";
      when 15006 => pixel <= "000000";
      when 15007 => pixel <= "000000";
      when 15008 => pixel <= "000000";
      when 15009 => pixel <= "000000";
      when 15010 => pixel <= "000000";
      when 15011 => pixel <= "000000";
      when 15012 => pixel <= "000000";
      when 15013 => pixel <= "000000";
      when 15014 => pixel <= "000000";
      when 15015 => pixel <= "000000";
      when 15016 => pixel <= "000000";
      when 15017 => pixel <= "000000";
      when 15018 => pixel <= "000000";
      when 15019 => pixel <= "000000";
      when 15020 => pixel <= "000000";
      when 15021 => pixel <= "000000";
      when 15022 => pixel <= "000000";
      when 15023 => pixel <= "000000";
      when 15024 => pixel <= "000000";
      when 15025 => pixel <= "000000";
      when 15026 => pixel <= "000000";
      when 15027 => pixel <= "000000";
      when 15028 => pixel <= "000000";
      when 15029 => pixel <= "000000";
      when 15030 => pixel <= "000000";
      when 15031 => pixel <= "000000";
      when 15032 => pixel <= "000000";
      when 15033 => pixel <= "000000";
      when 15034 => pixel <= "000000";
      when 15035 => pixel <= "000000";
      when 15036 => pixel <= "000000";
      when 15037 => pixel <= "000000";
      when 15038 => pixel <= "000000";
      when 15039 => pixel <= "000000";
      when 15040 => pixel <= "000000";
      when 15041 => pixel <= "000000";
      when 15042 => pixel <= "000000";
      when 15043 => pixel <= "000000";
      when 15044 => pixel <= "000000";
      when 15045 => pixel <= "000000";
      when 15046 => pixel <= "000000";
      when 15047 => pixel <= "000000";
      when 15048 => pixel <= "000000";
      when 15049 => pixel <= "000000";
      when 15050 => pixel <= "000000";
      when 15051 => pixel <= "000000";
      when 15052 => pixel <= "000000";
      when 15053 => pixel <= "000000";
      when 15054 => pixel <= "000000";
      when 15055 => pixel <= "000000";
      when 15056 => pixel <= "000000";
      when 15057 => pixel <= "000000";
      when 15058 => pixel <= "000000";
      when 15059 => pixel <= "000000";
      when 15060 => pixel <= "000000";
      when 15061 => pixel <= "000000";
      when 15062 => pixel <= "000000";
      when 15063 => pixel <= "000000";
      when 15064 => pixel <= "000000";
      when 15065 => pixel <= "000000";
      when 15066 => pixel <= "000000";
      when 15067 => pixel <= "000000";
      when 15068 => pixel <= "000000";
      when 15069 => pixel <= "000000";
      when 15070 => pixel <= "000000";
      when 15071 => pixel <= "000000";
      when 15072 => pixel <= "000000";
      when 15073 => pixel <= "000000";
      when 15074 => pixel <= "000000";
      when 15075 => pixel <= "000000";
      when 15076 => pixel <= "000000";
      when 15077 => pixel <= "000000";
      when 15078 => pixel <= "000000";
      when 15079 => pixel <= "000000";
      when 15080 => pixel <= "000000";
      when 15081 => pixel <= "000000";
      when 15082 => pixel <= "000000";
      when 15083 => pixel <= "000000";
      when 15084 => pixel <= "000000";
      when 15085 => pixel <= "000000";
      when 15086 => pixel <= "000000";
      when 15087 => pixel <= "000000";
      when 15088 => pixel <= "000000";
      when 15089 => pixel <= "000000";
      when 15090 => pixel <= "000000";
      when 15091 => pixel <= "000000";
      when 15092 => pixel <= "000000";
      when 15093 => pixel <= "000000";
      when 15094 => pixel <= "000000";
      when 15095 => pixel <= "000000";
      when 15096 => pixel <= "000000";
      when 15097 => pixel <= "000000";
      when 15098 => pixel <= "000000";
      when 15099 => pixel <= "000000";
      when 15100 => pixel <= "000000";
      when 15101 => pixel <= "000000";
      when 15102 => pixel <= "000000";
      when 15103 => pixel <= "000000";
      when 15104 => pixel <= "000000";
      when 15105 => pixel <= "000000";
      when 15106 => pixel <= "000000";
      when 15107 => pixel <= "000000";
      when 15108 => pixel <= "000000";
      when 15109 => pixel <= "000000";
      when 15110 => pixel <= "000000";
      when 15111 => pixel <= "000000";
      when 15112 => pixel <= "000000";
      when 15113 => pixel <= "000000";
      when 15114 => pixel <= "000000";
      when 15115 => pixel <= "000000";
      when 15116 => pixel <= "000000";
      when 15117 => pixel <= "000000";
      when 15118 => pixel <= "000000";
      when 15119 => pixel <= "000000";
      when 15120 => pixel <= "000000";
      when 15121 => pixel <= "000000";
      when 15122 => pixel <= "000000";
      when 15123 => pixel <= "000000";
      when 15124 => pixel <= "000000";
      when 15125 => pixel <= "000000";
      when 15126 => pixel <= "000000";
      when 15127 => pixel <= "000000";
      when 15128 => pixel <= "000000";
      when 15129 => pixel <= "000000";
      when 15130 => pixel <= "000000";
      when 15131 => pixel <= "000000";
      when 15132 => pixel <= "000000";
      when 15133 => pixel <= "000000";
      when 15134 => pixel <= "000000";
      when 15135 => pixel <= "000000";
      when 15136 => pixel <= "000000";
      when 15137 => pixel <= "000000";
      when 15138 => pixel <= "000000";
      when 15139 => pixel <= "000000";
      when 15140 => pixel <= "000000";
      when 15141 => pixel <= "000000";
      when 15142 => pixel <= "000000";
      when 15143 => pixel <= "000000";
      when 15144 => pixel <= "000000";
      when 15145 => pixel <= "000000";
      when 15146 => pixel <= "000000";
      when 15147 => pixel <= "000000";
      when 15148 => pixel <= "000000";
      when 15149 => pixel <= "000000";
      when 15150 => pixel <= "000000";
      when 15151 => pixel <= "000000";
      when 15152 => pixel <= "000000";
      when 15153 => pixel <= "000000";
      when 15154 => pixel <= "000000";
      when 15155 => pixel <= "000000";
      when 15156 => pixel <= "000000";
      when 15157 => pixel <= "000000";
      when 15158 => pixel <= "000000";
      when 15159 => pixel <= "000000";
      when 15160 => pixel <= "000000";
      when 15161 => pixel <= "000000";
      when 15162 => pixel <= "000000";
      when 15163 => pixel <= "000000";
      when 15164 => pixel <= "000000";
      when 15165 => pixel <= "000000";
      when 15166 => pixel <= "000000";
      when 15167 => pixel <= "000000";
      when 15168 => pixel <= "000000";
      when 15169 => pixel <= "000000";
      when 15170 => pixel <= "000000";
      when 15171 => pixel <= "000000";
      when 15172 => pixel <= "000000";
      when 15173 => pixel <= "000000";
      when 15174 => pixel <= "000000";
      when 15175 => pixel <= "000000";
      when 15176 => pixel <= "000000";
      when 15177 => pixel <= "000000";
      when 15178 => pixel <= "000000";
      when 15179 => pixel <= "000000";
      when 15180 => pixel <= "000000";
      when 15181 => pixel <= "000000";
      when 15182 => pixel <= "000000";
      when 15183 => pixel <= "000000";
      when 15184 => pixel <= "000000";
      when 15185 => pixel <= "000000";
      when 15186 => pixel <= "000000";
      when 15187 => pixel <= "000000";
      when 15188 => pixel <= "000000";
      when 15189 => pixel <= "000000";
      when 15190 => pixel <= "000000";
      when 15191 => pixel <= "000000";
      when 15192 => pixel <= "000000";
      when 15193 => pixel <= "000000";
      when 15194 => pixel <= "000000";
      when 15195 => pixel <= "000000";
      when 15196 => pixel <= "000000";
      when 15197 => pixel <= "000000";
      when 15198 => pixel <= "000000";
      when 15199 => pixel <= "000000";
      when 15200 => pixel <= "000000";
      when 15201 => pixel <= "000000";
      when 15202 => pixel <= "000000";
      when 15203 => pixel <= "000000";
      when 15204 => pixel <= "000000";
      when 15205 => pixel <= "000000";
      when 15206 => pixel <= "000000";
      when 15207 => pixel <= "000000";
      when 15208 => pixel <= "000000";
      when 15209 => pixel <= "000000";
      when 15210 => pixel <= "000000";
      when 15211 => pixel <= "000000";
      when 15212 => pixel <= "000000";
      when 15213 => pixel <= "000000";
      when 15214 => pixel <= "000000";
      when 15215 => pixel <= "000000";
      when 15216 => pixel <= "000000";
      when 15217 => pixel <= "000000";
      when 15218 => pixel <= "000000";
      when 15219 => pixel <= "000000";
      when 15220 => pixel <= "000000";
      when 15221 => pixel <= "000000";
      when 15222 => pixel <= "000000";
      when 15223 => pixel <= "000000";
      when 15224 => pixel <= "000000";
      when 15225 => pixel <= "000000";
      when 15226 => pixel <= "000000";
      when 15227 => pixel <= "000000";
      when 15228 => pixel <= "000000";
      when 15229 => pixel <= "000000";
      when 15230 => pixel <= "000000";
      when 15231 => pixel <= "000000";
      when 15232 => pixel <= "000000";
      when 15233 => pixel <= "000000";
      when 15234 => pixel <= "000000";
      when 15235 => pixel <= "000000";
      when 15236 => pixel <= "000000";
      when 15237 => pixel <= "000000";
      when 15238 => pixel <= "000000";
      when 15239 => pixel <= "000000";
      when 15240 => pixel <= "000000";
      when 15241 => pixel <= "000000";
      when 15242 => pixel <= "000000";
      when 15243 => pixel <= "000000";
      when 15244 => pixel <= "000000";
      when 15245 => pixel <= "000000";
      when 15246 => pixel <= "000000";
      when 15247 => pixel <= "000000";
      when 15248 => pixel <= "000000";
      when 15249 => pixel <= "000000";
      when 15250 => pixel <= "000000";
      when 15251 => pixel <= "000000";
      when 15252 => pixel <= "000000";
      when 15253 => pixel <= "000000";
      when 15254 => pixel <= "000000";
      when 15255 => pixel <= "000000";
      when 15256 => pixel <= "000000";
      when 15257 => pixel <= "000000";
      when 15258 => pixel <= "000000";
      when 15259 => pixel <= "000000";
      when 15260 => pixel <= "000000";
      when 15261 => pixel <= "000000";
      when 15262 => pixel <= "000000";
      when 15263 => pixel <= "000000";
      when 15264 => pixel <= "000000";
      when 15265 => pixel <= "000000";
      when 15266 => pixel <= "000000";
      when 15267 => pixel <= "000000";
      when 15268 => pixel <= "000000";
      when 15269 => pixel <= "000000";
      when 15270 => pixel <= "000000";
      when 15271 => pixel <= "000000";
      when 15272 => pixel <= "000000";
      when 15273 => pixel <= "000000";
      when 15274 => pixel <= "000000";
      when 15275 => pixel <= "000000";
      when 15276 => pixel <= "000000";
      when 15277 => pixel <= "000000";
      when 15278 => pixel <= "000000";
      when 15279 => pixel <= "000000";
      when 15280 => pixel <= "000000";
      when 15281 => pixel <= "000000";
      when 15282 => pixel <= "000000";
      when 15283 => pixel <= "000000";
      when 15284 => pixel <= "000000";
      when 15285 => pixel <= "000000";
      when 15286 => pixel <= "000000";
      when 15287 => pixel <= "000000";
      when 15288 => pixel <= "000000";
      when 15289 => pixel <= "000000";
      when 15290 => pixel <= "000000";
      when 15291 => pixel <= "000000";
      when 15292 => pixel <= "000000";
      when 15293 => pixel <= "000000";
      when 15294 => pixel <= "000000";
      when 15295 => pixel <= "000000";
      when 15296 => pixel <= "000000";
      when 15297 => pixel <= "000000";
      when 15298 => pixel <= "000000";
      when 15299 => pixel <= "000000";
      when 15300 => pixel <= "000000";
      when 15301 => pixel <= "000000";
      when 15302 => pixel <= "000000";
      when 15303 => pixel <= "000000";
      when 15304 => pixel <= "000000";
      when 15305 => pixel <= "000000";
      when 15306 => pixel <= "000000";
      when 15307 => pixel <= "000000";
      when 15308 => pixel <= "000000";
      when 15309 => pixel <= "000000";
      when 15310 => pixel <= "000000";
      when 15311 => pixel <= "000000";
      when 15312 => pixel <= "000000";
      when 15313 => pixel <= "000000";
      when 15314 => pixel <= "000000";
      when 15315 => pixel <= "000000";
      when 15316 => pixel <= "000000";
      when 15317 => pixel <= "000000";
      when 15318 => pixel <= "000000";
      when 15319 => pixel <= "000000";
      when 15320 => pixel <= "000000";
      when 15321 => pixel <= "000000";
      when 15322 => pixel <= "000000";
      when 15323 => pixel <= "000000";
      when 15324 => pixel <= "000000";
      when 15325 => pixel <= "000000";
      when 15326 => pixel <= "000000";
      when 15327 => pixel <= "000000";
      when 15328 => pixel <= "000000";
      when 15329 => pixel <= "000000";
      when 15330 => pixel <= "000000";
      when 15331 => pixel <= "000000";
      when 15332 => pixel <= "000000";
      when 15333 => pixel <= "000000";
      when 15334 => pixel <= "000000";
      when 15335 => pixel <= "000000";
      when 15336 => pixel <= "000000";
      when 15337 => pixel <= "000000";
      when 15338 => pixel <= "000000";
      when 15339 => pixel <= "000000";
      when 15340 => pixel <= "000000";
      when 15341 => pixel <= "000000";
      when 15342 => pixel <= "000000";
      when 15343 => pixel <= "000000";
      when 15344 => pixel <= "000000";
      when 15345 => pixel <= "000000";
      when 15346 => pixel <= "000000";
      when 15347 => pixel <= "000000";
      when 15348 => pixel <= "000000";
      when 15349 => pixel <= "000000";
      when 15350 => pixel <= "000000";
      when 15351 => pixel <= "000000";
      when 15352 => pixel <= "000000";
      when 15353 => pixel <= "000000";
      when 15354 => pixel <= "000000";
      when 15355 => pixel <= "000000";
      when 15356 => pixel <= "000000";
      when 15357 => pixel <= "000000";
      when 15358 => pixel <= "000000";
      when 15359 => pixel <= "000000";
      when 15360 => pixel <= "000000";
      when 15361 => pixel <= "000000";
      when 15362 => pixel <= "000000";
      when 15363 => pixel <= "000000";
      when 15364 => pixel <= "000000";
      when 15365 => pixel <= "000000";
      when 15366 => pixel <= "000000";
      when 15367 => pixel <= "000000";
      when 15368 => pixel <= "000000";
      when 15369 => pixel <= "000000";
      when 15370 => pixel <= "000000";
      when 15371 => pixel <= "000000";
      when 15372 => pixel <= "000000";
      when 15373 => pixel <= "000000";
      when 15374 => pixel <= "000000";
      when 15375 => pixel <= "000000";
      when 15376 => pixel <= "000000";
      when 15377 => pixel <= "000000";
      when 15378 => pixel <= "000000";
      when 15379 => pixel <= "000000";
      when 15380 => pixel <= "000000";
      when 15381 => pixel <= "000000";
      when 15382 => pixel <= "000000";
      when 15383 => pixel <= "000000";
      when 15384 => pixel <= "000000";
      when 15385 => pixel <= "000000";
      when 15386 => pixel <= "000000";
      when 15387 => pixel <= "000000";
      when 15388 => pixel <= "000000";
      when 15389 => pixel <= "000000";
      when 15390 => pixel <= "000000";
      when 15391 => pixel <= "000000";
      when 15392 => pixel <= "000000";
      when 15393 => pixel <= "000000";
      when 15394 => pixel <= "000000";
      when 15395 => pixel <= "000000";
      when 15396 => pixel <= "000000";
      when 15397 => pixel <= "000000";
      when 15398 => pixel <= "000000";
      when 15399 => pixel <= "000000";
      when 15400 => pixel <= "000000";
      when 15401 => pixel <= "000000";
      when 15402 => pixel <= "000000";
      when 15403 => pixel <= "000000";
      when 15404 => pixel <= "000000";
      when 15405 => pixel <= "000000";
      when 15406 => pixel <= "000000";
      when 15407 => pixel <= "000000";
      when 15408 => pixel <= "000000";
      when 15409 => pixel <= "000000";
      when 15410 => pixel <= "000000";
      when 15411 => pixel <= "000000";
      when 15412 => pixel <= "000000";
      when 15413 => pixel <= "000000";
      when 15414 => pixel <= "000000";
      when 15415 => pixel <= "000000";
      when 15416 => pixel <= "000000";
      when 15417 => pixel <= "000000";
      when 15418 => pixel <= "000000";
      when 15419 => pixel <= "000000";
      when 15420 => pixel <= "000000";
      when 15421 => pixel <= "000000";
      when 15422 => pixel <= "000000";
      when 15423 => pixel <= "000000";
      when 15424 => pixel <= "000000";
      when 15425 => pixel <= "000000";
      when 15426 => pixel <= "000000";
      when 15427 => pixel <= "000000";
      when 15428 => pixel <= "000000";
      when 15429 => pixel <= "000000";
      when 15430 => pixel <= "000000";
      when 15431 => pixel <= "000000";
      when 15432 => pixel <= "000000";
      when 15433 => pixel <= "000000";
      when 15434 => pixel <= "000000";
      when 15435 => pixel <= "000000";
      when 15436 => pixel <= "000000";
      when 15437 => pixel <= "000000";
      when 15438 => pixel <= "000000";
      when 15439 => pixel <= "000000";
      when 15440 => pixel <= "000000";
      when 15441 => pixel <= "000000";
      when 15442 => pixel <= "000000";
      when 15443 => pixel <= "000000";
      when 15444 => pixel <= "000000";
      when 15445 => pixel <= "000000";
      when 15446 => pixel <= "000000";
      when 15447 => pixel <= "000000";
      when 15448 => pixel <= "000000";
      when 15449 => pixel <= "000000";
      when 15450 => pixel <= "000000";
      when 15451 => pixel <= "000000";
      when 15452 => pixel <= "000000";
      when 15453 => pixel <= "000000";
      when 15454 => pixel <= "000000";
      when 15455 => pixel <= "000000";
      when 15456 => pixel <= "000000";
      when 15457 => pixel <= "000000";
      when 15458 => pixel <= "000000";
      when 15459 => pixel <= "000000";
      when 15460 => pixel <= "000000";
      when 15461 => pixel <= "000000";
      when 15462 => pixel <= "000000";
      when 15463 => pixel <= "000000";
      when 15464 => pixel <= "000000";
      when 15465 => pixel <= "000000";
      when 15466 => pixel <= "000000";
      when 15467 => pixel <= "000000";
      when 15468 => pixel <= "000000";
      when 15469 => pixel <= "000000";
      when 15470 => pixel <= "000000";
      when 15471 => pixel <= "000000";
      when 15472 => pixel <= "000000";
      when 15473 => pixel <= "000000";
      when 15474 => pixel <= "000000";
      when 15475 => pixel <= "000000";
      when 15476 => pixel <= "000000";
      when 15477 => pixel <= "000000";
      when 15478 => pixel <= "000000";
      when 15479 => pixel <= "000000";
      when 15480 => pixel <= "000000";
      when 15481 => pixel <= "000000";
      when 15482 => pixel <= "000000";
      when 15483 => pixel <= "000000";
      when 15484 => pixel <= "000000";
      when 15485 => pixel <= "000000";
      when 15486 => pixel <= "000000";
      when 15487 => pixel <= "000000";
      when 15488 => pixel <= "000000";
      when 15489 => pixel <= "000000";
      when 15490 => pixel <= "000000";
      when 15491 => pixel <= "000000";
      when 15492 => pixel <= "000000";
      when 15493 => pixel <= "000000";
      when 15494 => pixel <= "000000";
      when 15495 => pixel <= "000000";
      when 15496 => pixel <= "000000";
      when 15497 => pixel <= "000000";
      when 15498 => pixel <= "000000";
      when 15499 => pixel <= "000000";
      when 15500 => pixel <= "000000";
      when 15501 => pixel <= "000000";
      when 15502 => pixel <= "000000";
      when 15503 => pixel <= "000000";
      when 15504 => pixel <= "000000";
      when 15505 => pixel <= "000000";
      when 15506 => pixel <= "000000";
      when 15507 => pixel <= "000000";
      when 15508 => pixel <= "000000";
      when 15509 => pixel <= "000000";
      when 15510 => pixel <= "000000";
      when 15511 => pixel <= "000000";
      when 15512 => pixel <= "000000";
      when 15513 => pixel <= "000000";
      when 15514 => pixel <= "000000";
      when 15515 => pixel <= "000000";
      when 15516 => pixel <= "000000";
      when 15517 => pixel <= "000000";
      when 15518 => pixel <= "000000";
      when 15519 => pixel <= "000000";
      when 15520 => pixel <= "000000";
      when 15521 => pixel <= "000000";
      when 15522 => pixel <= "000000";
      when 15523 => pixel <= "000000";
      when 15524 => pixel <= "000000";
      when 15525 => pixel <= "000000";
      when 15526 => pixel <= "000000";
      when 15527 => pixel <= "000000";
      when 15528 => pixel <= "000000";
      when 15529 => pixel <= "000000";
      when 15530 => pixel <= "000000";
      when 15531 => pixel <= "000000";
      when 15532 => pixel <= "000000";
      when 15533 => pixel <= "000000";
      when 15534 => pixel <= "000000";
      when 15535 => pixel <= "000000";
      when 15536 => pixel <= "000000";
      when 15537 => pixel <= "000000";
      when 15538 => pixel <= "000000";
      when 15539 => pixel <= "000000";
      when 15540 => pixel <= "000000";
      when 15541 => pixel <= "000000";
      when 15542 => pixel <= "000000";
      when 15543 => pixel <= "000000";
      when 15544 => pixel <= "000000";
      when 15545 => pixel <= "000000";
      when 15546 => pixel <= "000000";
      when 15547 => pixel <= "000000";
      when 15548 => pixel <= "000000";
      when 15549 => pixel <= "000000";
      when 15550 => pixel <= "000000";
      when 15551 => pixel <= "000000";
      when 15552 => pixel <= "000000";
      when 15553 => pixel <= "000000";
      when 15554 => pixel <= "000000";
      when 15555 => pixel <= "000000";
      when 15556 => pixel <= "000000";
      when 15557 => pixel <= "000000";
      when 15558 => pixel <= "000000";
      when 15559 => pixel <= "000000";
      when 15560 => pixel <= "000000";
      when 15561 => pixel <= "000000";
      when 15562 => pixel <= "000000";
      when 15563 => pixel <= "000000";
      when 15564 => pixel <= "000000";
      when 15565 => pixel <= "000000";
      when 15566 => pixel <= "000000";
      when 15567 => pixel <= "000000";
      when 15568 => pixel <= "000000";
      when 15569 => pixel <= "000000";
      when 15570 => pixel <= "000000";
      when 15571 => pixel <= "000000";
      when 15572 => pixel <= "000000";
      when 15573 => pixel <= "000000";
      when 15574 => pixel <= "000000";
      when 15575 => pixel <= "000000";
      when 15576 => pixel <= "000000";
      when 15577 => pixel <= "000000";
      when 15578 => pixel <= "000000";
      when 15579 => pixel <= "000000";
      when 15580 => pixel <= "000000";
      when 15581 => pixel <= "000000";
      when 15582 => pixel <= "000000";
      when 15583 => pixel <= "000000";
      when 15584 => pixel <= "000000";
      when 15585 => pixel <= "000000";
      when 15586 => pixel <= "000000";
      when 15587 => pixel <= "000000";
      when 15588 => pixel <= "000000";
      when 15589 => pixel <= "000000";
      when 15590 => pixel <= "000000";
      when 15591 => pixel <= "000000";
      when 15592 => pixel <= "000000";
      when 15593 => pixel <= "000000";
      when 15594 => pixel <= "000000";
      when 15595 => pixel <= "000000";
      when 15596 => pixel <= "000000";
      when 15597 => pixel <= "000000";
      when 15598 => pixel <= "000000";
      when 15599 => pixel <= "000000";
      when 15600 => pixel <= "000000";
      when 15601 => pixel <= "000000";
      when 15602 => pixel <= "000000";
      when 15603 => pixel <= "000000";
      when 15604 => pixel <= "000000";
      when 15605 => pixel <= "000000";
      when 15606 => pixel <= "000000";
      when 15607 => pixel <= "000000";
      when 15608 => pixel <= "000000";
      when 15609 => pixel <= "000000";
      when 15610 => pixel <= "000000";
      when 15611 => pixel <= "000000";
      when 15612 => pixel <= "000000";
      when 15613 => pixel <= "000000";
      when 15614 => pixel <= "000000";
      when 15615 => pixel <= "000000";
      when 15616 => pixel <= "000000";
      when 15617 => pixel <= "000000";
      when 15618 => pixel <= "000000";
      when 15619 => pixel <= "000000";
      when 15620 => pixel <= "000000";
      when 15621 => pixel <= "000000";
      when 15622 => pixel <= "000000";
      when 15623 => pixel <= "000000";
      when 15624 => pixel <= "000000";
      when 15625 => pixel <= "000000";
      when 15626 => pixel <= "000000";
      when 15627 => pixel <= "000000";
      when 15628 => pixel <= "000000";
      when 15629 => pixel <= "000000";
      when 15630 => pixel <= "000000";
      when 15631 => pixel <= "000000";
      when 15632 => pixel <= "000000";
      when 15633 => pixel <= "000000";
      when 15634 => pixel <= "000000";
      when 15635 => pixel <= "000000";
      when 15636 => pixel <= "000000";
      when 15637 => pixel <= "000000";
      when 15638 => pixel <= "000000";
      when 15639 => pixel <= "000000";
      when 15640 => pixel <= "000000";
      when 15641 => pixel <= "000000";
      when 15642 => pixel <= "000000";
      when 15643 => pixel <= "000000";
      when 15644 => pixel <= "000000";
      when 15645 => pixel <= "000000";
      when 15646 => pixel <= "000000";
      when 15647 => pixel <= "000000";
      when 15648 => pixel <= "000000";
      when 15649 => pixel <= "000000";
      when 15650 => pixel <= "000000";
      when 15651 => pixel <= "000000";
      when 15652 => pixel <= "000000";
      when 15653 => pixel <= "000000";
      when 15654 => pixel <= "000000";
      when 15655 => pixel <= "000000";
      when 15656 => pixel <= "000000";
      when 15657 => pixel <= "000000";
      when 15658 => pixel <= "000000";
      when 15659 => pixel <= "000000";
      when 15660 => pixel <= "000000";
      when 15661 => pixel <= "000000";
      when 15662 => pixel <= "000000";
      when 15663 => pixel <= "000000";
      when 15664 => pixel <= "000000";
      when 15665 => pixel <= "000000";
      when 15666 => pixel <= "000000";
      when 15667 => pixel <= "000000";
      when 15668 => pixel <= "000000";
      when 15669 => pixel <= "000000";
      when 15670 => pixel <= "000000";
      when 15671 => pixel <= "000000";
      when 15672 => pixel <= "000000";
      when 15673 => pixel <= "000000";
      when 15674 => pixel <= "000000";
      when 15675 => pixel <= "000000";
      when 15676 => pixel <= "000000";
      when 15677 => pixel <= "000000";
      when 15678 => pixel <= "000000";
      when 15679 => pixel <= "000000";
      when 15680 => pixel <= "000000";
      when 15681 => pixel <= "000000";
      when 15682 => pixel <= "000000";
      when 15683 => pixel <= "000000";
      when 15684 => pixel <= "000000";
      when 15685 => pixel <= "000000";
      when 15686 => pixel <= "000000";
      when 15687 => pixel <= "000000";
      when 15688 => pixel <= "000000";
      when 15689 => pixel <= "000000";
      when 15690 => pixel <= "000000";
      when 15691 => pixel <= "000000";
      when 15692 => pixel <= "000000";
      when 15693 => pixel <= "000000";
      when 15694 => pixel <= "000000";
      when 15695 => pixel <= "000000";
      when 15696 => pixel <= "000000";
      when 15697 => pixel <= "000000";
      when 15698 => pixel <= "000000";
      when 15699 => pixel <= "000000";
      when 15700 => pixel <= "000000";
      when 15701 => pixel <= "000000";
      when 15702 => pixel <= "000000";
      when 15703 => pixel <= "000000";
      when 15704 => pixel <= "000000";
      when 15705 => pixel <= "000000";
      when 15706 => pixel <= "000000";
      when 15707 => pixel <= "000000";
      when 15708 => pixel <= "000000";
      when 15709 => pixel <= "000000";
      when 15710 => pixel <= "000000";
      when 15711 => pixel <= "000000";
      when 15712 => pixel <= "000000";
      when 15713 => pixel <= "000000";
      when 15714 => pixel <= "000000";
      when 15715 => pixel <= "000000";
      when 15716 => pixel <= "000000";
      when 15717 => pixel <= "000000";
      when 15718 => pixel <= "000000";
      when 15719 => pixel <= "000000";
      when 15720 => pixel <= "000000";
      when 15721 => pixel <= "000000";
      when 15722 => pixel <= "000000";
      when 15723 => pixel <= "000000";
      when 15724 => pixel <= "000000";
      when 15725 => pixel <= "000000";
      when 15726 => pixel <= "000000";
      when 15727 => pixel <= "000000";
      when 15728 => pixel <= "000000";
      when 15729 => pixel <= "000000";
      when 15730 => pixel <= "000000";
      when 15731 => pixel <= "000000";
      when 15732 => pixel <= "000000";
      when 15733 => pixel <= "000000";
      when 15734 => pixel <= "000000";
      when 15735 => pixel <= "000000";
      when 15736 => pixel <= "000000";
      when 15737 => pixel <= "000000";
      when 15738 => pixel <= "000000";
      when 15739 => pixel <= "000000";
      when 15740 => pixel <= "000000";
      when 15741 => pixel <= "000000";
      when 15742 => pixel <= "000000";
      when 15743 => pixel <= "000000";
      when 15744 => pixel <= "000000";
      when 15745 => pixel <= "000000";
      when 15746 => pixel <= "000000";
      when 15747 => pixel <= "000000";
      when 15748 => pixel <= "000000";
      when 15749 => pixel <= "000000";
      when 15750 => pixel <= "000000";
      when 15751 => pixel <= "000000";
      when 15752 => pixel <= "000000";
      when 15753 => pixel <= "000000";
      when 15754 => pixel <= "000000";
      when 15755 => pixel <= "000000";
      when 15756 => pixel <= "000000";
      when 15757 => pixel <= "000000";
      when 15758 => pixel <= "000000";
      when 15759 => pixel <= "000000";
      when 15760 => pixel <= "000000";
      when 15761 => pixel <= "000000";
      when 15762 => pixel <= "000000";
      when 15763 => pixel <= "000000";
      when 15764 => pixel <= "000000";
      when 15765 => pixel <= "000000";
      when 15766 => pixel <= "000000";
      when 15767 => pixel <= "000000";
      when 15768 => pixel <= "000000";
      when 15769 => pixel <= "000000";
      when 15770 => pixel <= "000000";
      when 15771 => pixel <= "000000";
      when 15772 => pixel <= "000000";
      when 15773 => pixel <= "000000";
      when 15774 => pixel <= "000000";
      when 15775 => pixel <= "000000";
      when 15776 => pixel <= "000000";
      when 15777 => pixel <= "000000";
      when 15778 => pixel <= "000000";
      when 15779 => pixel <= "000000";
      when 15780 => pixel <= "000000";
      when 15781 => pixel <= "000000";
      when 15782 => pixel <= "000000";
      when 15783 => pixel <= "000000";
      when 15784 => pixel <= "000000";
      when 15785 => pixel <= "000000";
      when 15786 => pixel <= "000000";
      when 15787 => pixel <= "000000";
      when 15788 => pixel <= "000000";
      when 15789 => pixel <= "000000";
      when 15790 => pixel <= "000000";
      when 15791 => pixel <= "000000";
      when 15792 => pixel <= "000000";
      when 15793 => pixel <= "000000";
      when 15794 => pixel <= "000000";
      when 15795 => pixel <= "000000";
      when 15796 => pixel <= "000000";
      when 15797 => pixel <= "000000";
      when 15798 => pixel <= "000000";
      when 15799 => pixel <= "000000";
      when 15800 => pixel <= "000000";
      when 15801 => pixel <= "000000";
      when 15802 => pixel <= "000000";
      when 15803 => pixel <= "000000";
      when 15804 => pixel <= "000000";
      when 15805 => pixel <= "000000";
      when 15806 => pixel <= "000000";
      when 15807 => pixel <= "000000";
      when 15808 => pixel <= "000000";
      when 15809 => pixel <= "000000";
      when 15810 => pixel <= "000000";
      when 15811 => pixel <= "000000";
      when 15812 => pixel <= "000000";
      when 15813 => pixel <= "000000";
      when 15814 => pixel <= "000000";
      when 15815 => pixel <= "000000";
      when 15816 => pixel <= "000000";
      when 15817 => pixel <= "000000";
      when 15818 => pixel <= "000000";
      when 15819 => pixel <= "000000";
      when 15820 => pixel <= "000000";
      when 15821 => pixel <= "000000";
      when 15822 => pixel <= "000000";
      when 15823 => pixel <= "000000";
      when 15824 => pixel <= "000000";
      when 15825 => pixel <= "000000";
      when 15826 => pixel <= "000000";
      when 15827 => pixel <= "000000";
      when 15828 => pixel <= "000000";
      when 15829 => pixel <= "000000";
      when 15830 => pixel <= "000000";
      when 15831 => pixel <= "000000";
      when 15832 => pixel <= "000000";
      when 15833 => pixel <= "000000";
      when 15834 => pixel <= "000000";
      when 15835 => pixel <= "000000";
      when 15836 => pixel <= "000000";
      when 15837 => pixel <= "000000";
      when 15838 => pixel <= "000000";
      when 15839 => pixel <= "000000";
      when 15840 => pixel <= "000000";
      when 15841 => pixel <= "000000";
      when 15842 => pixel <= "000000";
      when 15843 => pixel <= "000000";
      when 15844 => pixel <= "000000";
      when 15845 => pixel <= "000000";
      when 15846 => pixel <= "000000";
      when 15847 => pixel <= "000000";
      when 15848 => pixel <= "000000";
      when 15849 => pixel <= "000000";
      when 15850 => pixel <= "000000";
      when 15851 => pixel <= "000000";
      when 15852 => pixel <= "000000";
      when 15853 => pixel <= "000000";
      when 15854 => pixel <= "000000";
      when 15855 => pixel <= "000000";
      when 15856 => pixel <= "000000";
      when 15857 => pixel <= "000000";
      when 15858 => pixel <= "000000";
      when 15859 => pixel <= "000000";
      when 15860 => pixel <= "000000";
      when 15861 => pixel <= "000000";
      when 15862 => pixel <= "000000";
      when 15863 => pixel <= "000000";
      when 15864 => pixel <= "000000";
      when 15865 => pixel <= "000000";
      when 15866 => pixel <= "000000";
      when 15867 => pixel <= "000000";
      when 15868 => pixel <= "000000";
      when 15869 => pixel <= "000000";
      when 15870 => pixel <= "000000";
      when 15871 => pixel <= "000000";
      when 15872 => pixel <= "000000";
      when 15873 => pixel <= "000000";
      when 15874 => pixel <= "000000";
      when 15875 => pixel <= "000000";
      when 15876 => pixel <= "000000";
      when 15877 => pixel <= "000000";
      when 15878 => pixel <= "000000";
      when 15879 => pixel <= "000000";
      when 15880 => pixel <= "000000";
      when 15881 => pixel <= "000000";
      when 15882 => pixel <= "000000";
      when 15883 => pixel <= "000000";
      when 15884 => pixel <= "000000";
      when 15885 => pixel <= "000000";
      when 15886 => pixel <= "000000";
      when 15887 => pixel <= "000000";
      when 15888 => pixel <= "000000";
      when 15889 => pixel <= "000000";
      when 15890 => pixel <= "000000";
      when 15891 => pixel <= "000000";
      when 15892 => pixel <= "000000";
      when 15893 => pixel <= "000000";
      when 15894 => pixel <= "000000";
      when 15895 => pixel <= "000000";
      when 15896 => pixel <= "000000";
      when 15897 => pixel <= "000000";
      when 15898 => pixel <= "000000";
      when 15899 => pixel <= "000000";
      when 15900 => pixel <= "000000";
      when 15901 => pixel <= "000000";
      when 15902 => pixel <= "000000";
      when 15903 => pixel <= "000000";
      when 15904 => pixel <= "000000";
      when 15905 => pixel <= "000000";
      when 15906 => pixel <= "000000";
      when 15907 => pixel <= "000000";
      when 15908 => pixel <= "000000";
      when 15909 => pixel <= "000000";
      when 15910 => pixel <= "000000";
      when 15911 => pixel <= "000000";
      when 15912 => pixel <= "000000";
      when 15913 => pixel <= "000000";
      when 15914 => pixel <= "000000";
      when 15915 => pixel <= "000000";
      when 15916 => pixel <= "000000";
      when 15917 => pixel <= "000000";
      when 15918 => pixel <= "000000";
      when 15919 => pixel <= "000000";
      when 15920 => pixel <= "000000";
      when 15921 => pixel <= "000000";
      when 15922 => pixel <= "000000";
      when 15923 => pixel <= "000000";
      when 15924 => pixel <= "000000";
      when 15925 => pixel <= "000000";
      when 15926 => pixel <= "000000";
      when 15927 => pixel <= "000000";
      when 15928 => pixel <= "000000";
      when 15929 => pixel <= "000000";
      when 15930 => pixel <= "000000";
      when 15931 => pixel <= "000000";
      when 15932 => pixel <= "000000";
      when 15933 => pixel <= "000000";
      when 15934 => pixel <= "000000";
      when 15935 => pixel <= "000000";
      when 15936 => pixel <= "000000";
      when 15937 => pixel <= "000000";
      when 15938 => pixel <= "000000";
      when 15939 => pixel <= "000000";
      when 15940 => pixel <= "000000";
      when 15941 => pixel <= "000000";
      when 15942 => pixel <= "000000";
      when 15943 => pixel <= "000000";
      when 15944 => pixel <= "000000";
      when 15945 => pixel <= "000000";
      when 15946 => pixel <= "000000";
      when 15947 => pixel <= "000000";
      when 15948 => pixel <= "000000";
      when 15949 => pixel <= "000000";
      when 15950 => pixel <= "000000";
      when 15951 => pixel <= "000000";
      when 15952 => pixel <= "000000";
      when 15953 => pixel <= "000000";
      when 15954 => pixel <= "000000";
      when 15955 => pixel <= "000000";
      when 15956 => pixel <= "000000";
      when 15957 => pixel <= "000000";
      when 15958 => pixel <= "000000";
      when 15959 => pixel <= "000000";
      when 15960 => pixel <= "000000";
      when 15961 => pixel <= "000000";
      when 15962 => pixel <= "000000";
      when 15963 => pixel <= "000000";
      when 15964 => pixel <= "000000";
      when 15965 => pixel <= "000000";
      when 15966 => pixel <= "000000";
      when 15967 => pixel <= "000000";
      when 15968 => pixel <= "000000";
      when 15969 => pixel <= "000000";
      when 15970 => pixel <= "000000";
      when 15971 => pixel <= "000000";
      when 15972 => pixel <= "000000";
      when 15973 => pixel <= "000000";
      when 15974 => pixel <= "000000";
      when 15975 => pixel <= "000000";
      when 15976 => pixel <= "000000";
      when 15977 => pixel <= "000000";
      when 15978 => pixel <= "000000";
      when 15979 => pixel <= "000000";
      when 15980 => pixel <= "000000";
      when 15981 => pixel <= "000000";
      when 15982 => pixel <= "000000";
      when 15983 => pixel <= "000000";
      when 15984 => pixel <= "000000";
      when 15985 => pixel <= "000000";
      when 15986 => pixel <= "000000";
      when 15987 => pixel <= "000000";
      when 15988 => pixel <= "000000";
      when 15989 => pixel <= "000000";
      when 15990 => pixel <= "000000";
      when 15991 => pixel <= "000000";
      when 15992 => pixel <= "000000";
      when 15993 => pixel <= "000000";
      when 15994 => pixel <= "000000";
      when 15995 => pixel <= "000000";
      when 15996 => pixel <= "000000";
      when 15997 => pixel <= "000000";
      when 15998 => pixel <= "000000";
      when 15999 => pixel <= "000000";
      when 16000 => pixel <= "000000";
      when 16001 => pixel <= "000000";
      when 16002 => pixel <= "000000";
      when 16003 => pixel <= "000000";
      when 16004 => pixel <= "000000";
      when 16005 => pixel <= "000000";
      when 16006 => pixel <= "000000";
      when 16007 => pixel <= "000000";
      when 16008 => pixel <= "000000";
      when 16009 => pixel <= "000000";
      when 16010 => pixel <= "000000";
      when 16011 => pixel <= "000000";
      when 16012 => pixel <= "000000";
      when 16013 => pixel <= "000000";
      when 16014 => pixel <= "000000";
      when 16015 => pixel <= "000000";
      when 16016 => pixel <= "000000";
      when 16017 => pixel <= "000000";
      when 16018 => pixel <= "000000";
      when 16019 => pixel <= "000000";
      when 16020 => pixel <= "000000";
      when 16021 => pixel <= "000000";
      when 16022 => pixel <= "000000";
      when 16023 => pixel <= "000000";
      when 16024 => pixel <= "000000";
      when 16025 => pixel <= "000000";
      when 16026 => pixel <= "000000";
      when 16027 => pixel <= "000000";
      when 16028 => pixel <= "000000";
      when 16029 => pixel <= "000000";
      when 16030 => pixel <= "000000";
      when 16031 => pixel <= "000000";
      when 16032 => pixel <= "000000";
      when 16033 => pixel <= "000000";
      when 16034 => pixel <= "000000";
      when 16035 => pixel <= "000000";
      when 16036 => pixel <= "000000";
      when 16037 => pixel <= "000000";
      when 16038 => pixel <= "000000";
      when 16039 => pixel <= "000000";
      when 16040 => pixel <= "000000";
      when 16041 => pixel <= "000000";
      when 16042 => pixel <= "000000";
      when 16043 => pixel <= "000000";
      when 16044 => pixel <= "000000";
      when 16045 => pixel <= "000000";
      when 16046 => pixel <= "000000";
      when 16047 => pixel <= "000000";
      when 16048 => pixel <= "000000";
      when 16049 => pixel <= "000000";
      when 16050 => pixel <= "000000";
      when 16051 => pixel <= "000000";
      when 16052 => pixel <= "000000";
      when 16053 => pixel <= "000000";
      when 16054 => pixel <= "000000";
      when 16055 => pixel <= "000000";
      when 16056 => pixel <= "000000";
      when 16057 => pixel <= "000000";
      when 16058 => pixel <= "000000";
      when 16059 => pixel <= "000000";
      when 16060 => pixel <= "000000";
      when 16061 => pixel <= "000000";
      when 16062 => pixel <= "000000";
      when 16063 => pixel <= "000000";
      when 16064 => pixel <= "000000";
      when 16065 => pixel <= "000000";
      when 16066 => pixel <= "000000";
      when 16067 => pixel <= "000000";
      when 16068 => pixel <= "000000";
      when 16069 => pixel <= "000000";
      when 16070 => pixel <= "000000";
      when 16071 => pixel <= "000000";
      when 16072 => pixel <= "000000";
      when 16073 => pixel <= "000000";
      when 16074 => pixel <= "000000";
      when 16075 => pixel <= "000000";
      when 16076 => pixel <= "000000";
      when 16077 => pixel <= "000000";
      when 16078 => pixel <= "000000";
      when 16079 => pixel <= "000000";
      when 16080 => pixel <= "000000";
      when 16081 => pixel <= "000000";
      when 16082 => pixel <= "000000";
      when 16083 => pixel <= "000000";
      when 16084 => pixel <= "000000";
      when 16085 => pixel <= "000000";
      when 16086 => pixel <= "000000";
      when 16087 => pixel <= "000000";
      when 16088 => pixel <= "000000";
      when 16089 => pixel <= "000000";
      when 16090 => pixel <= "000000";
      when 16091 => pixel <= "000000";
      when 16092 => pixel <= "000000";
      when 16093 => pixel <= "000000";
      when 16094 => pixel <= "000000";
      when 16095 => pixel <= "000000";
      when 16096 => pixel <= "000000";
      when 16097 => pixel <= "000000";
      when 16098 => pixel <= "000000";
      when 16099 => pixel <= "000000";
      when 16100 => pixel <= "000000";
      when 16101 => pixel <= "000000";
      when 16102 => pixel <= "000000";
      when 16103 => pixel <= "000000";
      when 16104 => pixel <= "000000";
      when 16105 => pixel <= "000000";
      when 16106 => pixel <= "000000";
      when 16107 => pixel <= "000000";
      when 16108 => pixel <= "000000";
      when 16109 => pixel <= "000000";
      when 16110 => pixel <= "000000";
      when 16111 => pixel <= "000000";
      when 16112 => pixel <= "000000";
      when 16113 => pixel <= "000000";
      when 16114 => pixel <= "000000";
      when 16115 => pixel <= "000000";
      when 16116 => pixel <= "000000";
      when 16117 => pixel <= "000000";
      when 16118 => pixel <= "000000";
      when 16119 => pixel <= "000000";
      when 16120 => pixel <= "000000";
      when 16121 => pixel <= "000000";
      when 16122 => pixel <= "000000";
      when 16123 => pixel <= "000000";
      when 16124 => pixel <= "000000";
      when 16125 => pixel <= "000000";
      when 16126 => pixel <= "000000";
      when 16127 => pixel <= "000000";
      when 16128 => pixel <= "000000";
      when 16129 => pixel <= "000000";
      when 16130 => pixel <= "000000";
      when 16131 => pixel <= "000000";
      when 16132 => pixel <= "000000";
      when 16133 => pixel <= "000000";
      when 16134 => pixel <= "000000";
      when 16135 => pixel <= "000000";
      when 16136 => pixel <= "000000";
      when 16137 => pixel <= "000000";
      when 16138 => pixel <= "000000";
      when 16139 => pixel <= "000000";
      when 16140 => pixel <= "000000";
      when 16141 => pixel <= "000000";
      when 16142 => pixel <= "000000";
      when 16143 => pixel <= "000000";
      when 16144 => pixel <= "000000";
      when 16145 => pixel <= "000000";
      when 16146 => pixel <= "000000";
      when 16147 => pixel <= "000000";
      when 16148 => pixel <= "000000";
      when 16149 => pixel <= "000000";
      when 16150 => pixel <= "000000";
      when 16151 => pixel <= "000000";
      when 16152 => pixel <= "000000";
      when 16153 => pixel <= "000000";
      when 16154 => pixel <= "000000";
      when 16155 => pixel <= "000000";
      when 16156 => pixel <= "000000";
      when 16157 => pixel <= "000000";
      when 16158 => pixel <= "000000";
      when 16159 => pixel <= "000000";
      when 16160 => pixel <= "000000";
      when 16161 => pixel <= "000000";
      when 16162 => pixel <= "000000";
      when 16163 => pixel <= "000000";
      when 16164 => pixel <= "000000";
      when 16165 => pixel <= "000000";
      when 16166 => pixel <= "000000";
      when 16167 => pixel <= "000000";
      when 16168 => pixel <= "000000";
      when 16169 => pixel <= "000000";
      when 16170 => pixel <= "000000";
      when 16171 => pixel <= "000000";
      when 16172 => pixel <= "000000";
      when 16173 => pixel <= "000000";
      when 16174 => pixel <= "000000";
      when 16175 => pixel <= "000000";
      when 16176 => pixel <= "000000";
      when 16177 => pixel <= "000000";
      when 16178 => pixel <= "000000";
      when 16179 => pixel <= "000000";
      when 16180 => pixel <= "000000";
      when 16181 => pixel <= "000000";
      when 16182 => pixel <= "000000";
      when 16183 => pixel <= "000000";
      when 16184 => pixel <= "000000";
      when 16185 => pixel <= "000000";
      when 16186 => pixel <= "000000";
      when 16187 => pixel <= "000000";
      when 16188 => pixel <= "000000";
      when 16189 => pixel <= "000000";
      when 16190 => pixel <= "000000";
      when 16191 => pixel <= "000000";
      when 16192 => pixel <= "000000";
      when 16193 => pixel <= "000000";
      when 16194 => pixel <= "000000";
      when 16195 => pixel <= "000000";
      when 16196 => pixel <= "000000";
      when 16197 => pixel <= "000000";
      when 16198 => pixel <= "000000";
      when 16199 => pixel <= "000000";
      when 16200 => pixel <= "000000";
      when 16201 => pixel <= "000000";
      when 16202 => pixel <= "000000";
      when 16203 => pixel <= "000000";
      when 16204 => pixel <= "000000";
      when 16205 => pixel <= "000000";
      when 16206 => pixel <= "000000";
      when 16207 => pixel <= "000000";
      when 16208 => pixel <= "000000";
      when 16209 => pixel <= "000000";
      when 16210 => pixel <= "000000";
      when 16211 => pixel <= "000000";
      when 16212 => pixel <= "000000";
      when 16213 => pixel <= "000000";
      when 16214 => pixel <= "000000";
      when 16215 => pixel <= "000000";
      when 16216 => pixel <= "000000";
      when 16217 => pixel <= "000000";
      when 16218 => pixel <= "000000";
      when 16219 => pixel <= "000000";
      when 16220 => pixel <= "000000";
      when 16221 => pixel <= "000000";
      when 16222 => pixel <= "000000";
      when 16223 => pixel <= "000000";
      when 16224 => pixel <= "000000";
      when 16225 => pixel <= "000000";
      when 16226 => pixel <= "000000";
      when 16227 => pixel <= "000000";
      when 16228 => pixel <= "000000";
      when 16229 => pixel <= "000000";
      when 16230 => pixel <= "000000";
      when 16231 => pixel <= "000000";
      when 16232 => pixel <= "000000";
      when 16233 => pixel <= "000000";
      when 16234 => pixel <= "000000";
      when 16235 => pixel <= "000000";
      when 16236 => pixel <= "000000";
      when 16237 => pixel <= "000000";
      when 16238 => pixel <= "000000";
      when 16239 => pixel <= "000000";
      when 16240 => pixel <= "000000";
      when 16241 => pixel <= "000000";
      when 16242 => pixel <= "000000";
      when 16243 => pixel <= "000000";
      when 16244 => pixel <= "000000";
      when 16245 => pixel <= "000000";
      when 16246 => pixel <= "000000";
      when 16247 => pixel <= "000000";
      when 16248 => pixel <= "000000";
      when 16249 => pixel <= "000000";
      when 16250 => pixel <= "000000";
      when 16251 => pixel <= "000000";
      when 16252 => pixel <= "000000";
      when 16253 => pixel <= "000000";
      when 16254 => pixel <= "000000";
      when 16255 => pixel <= "000000";
      when 16256 => pixel <= "000000";
      when 16257 => pixel <= "000000";
      when 16258 => pixel <= "000000";
      when 16259 => pixel <= "000000";
      when 16260 => pixel <= "000000";
      when 16261 => pixel <= "000000";
      when 16262 => pixel <= "000000";
      when 16263 => pixel <= "000000";
      when 16264 => pixel <= "000000";
      when 16265 => pixel <= "000000";
      when 16266 => pixel <= "000000";
      when 16267 => pixel <= "000000";
      when 16268 => pixel <= "000000";
      when 16269 => pixel <= "000000";
      when 16270 => pixel <= "000000";
      when 16271 => pixel <= "000000";
      when 16272 => pixel <= "000000";
      when 16273 => pixel <= "000000";
      when 16274 => pixel <= "000000";
      when 16275 => pixel <= "000000";
      when 16276 => pixel <= "000000";
      when 16277 => pixel <= "000000";
      when 16278 => pixel <= "000000";
      when 16279 => pixel <= "000000";
      when 16280 => pixel <= "000000";
      when 16281 => pixel <= "000000";
      when 16282 => pixel <= "000000";
      when 16283 => pixel <= "000000";
      when 16284 => pixel <= "000000";
      when 16285 => pixel <= "000000";
      when 16286 => pixel <= "000000";
      when 16287 => pixel <= "000000";
      when 16288 => pixel <= "000000";
      when 16289 => pixel <= "000000";
      when 16290 => pixel <= "000000";
      when 16291 => pixel <= "000000";
      when 16292 => pixel <= "000000";
      when 16293 => pixel <= "000000";
      when 16294 => pixel <= "000000";
      when 16295 => pixel <= "000000";
      when 16296 => pixel <= "000000";
      when 16297 => pixel <= "000000";
      when 16298 => pixel <= "000000";
      when 16299 => pixel <= "000000";
      when 16300 => pixel <= "000000";
      when 16301 => pixel <= "000000";
      when 16302 => pixel <= "000000";
      when 16303 => pixel <= "000000";
      when 16304 => pixel <= "000000";
      when 16305 => pixel <= "000000";
      when 16306 => pixel <= "000000";
      when 16307 => pixel <= "000000";
      when 16308 => pixel <= "000000";
      when 16309 => pixel <= "000000";
      when 16310 => pixel <= "000000";
      when 16311 => pixel <= "000000";
      when 16312 => pixel <= "000000";
      when 16313 => pixel <= "000000";
      when 16314 => pixel <= "000000";
      when 16315 => pixel <= "000000";
      when 16316 => pixel <= "000000";
      when 16317 => pixel <= "000000";
      when 16318 => pixel <= "000000";
      when 16319 => pixel <= "000000";
      when 16320 => pixel <= "000000";
      when 16321 => pixel <= "000000";
      when 16322 => pixel <= "000000";
      when 16323 => pixel <= "000000";
      when 16324 => pixel <= "000000";
      when 16325 => pixel <= "000000";
      when 16326 => pixel <= "000000";
      when 16327 => pixel <= "000000";
      when 16328 => pixel <= "000000";
      when 16329 => pixel <= "000000";
      when 16330 => pixel <= "000000";
      when 16331 => pixel <= "000000";
      when 16332 => pixel <= "000000";
      when 16333 => pixel <= "000000";
      when 16334 => pixel <= "000000";
      when 16335 => pixel <= "000000";
      when 16336 => pixel <= "000000";
      when 16337 => pixel <= "000000";
      when 16338 => pixel <= "000000";
      when 16339 => pixel <= "000000";
      when 16340 => pixel <= "000000";
      when 16341 => pixel <= "000000";
      when 16342 => pixel <= "000000";
      when 16343 => pixel <= "000000";
      when 16344 => pixel <= "000000";
      when 16345 => pixel <= "000000";
      when 16346 => pixel <= "000000";
      when 16347 => pixel <= "000000";
      when 16348 => pixel <= "000000";
      when 16349 => pixel <= "000000";
      when 16350 => pixel <= "000000";
      when 16351 => pixel <= "000000";
      when 16352 => pixel <= "000000";
      when 16353 => pixel <= "000000";
      when 16354 => pixel <= "000000";
      when 16355 => pixel <= "000000";
      when 16356 => pixel <= "000000";
      when 16357 => pixel <= "000000";
      when 16358 => pixel <= "000000";
      when 16359 => pixel <= "000000";
      when 16360 => pixel <= "000000";
      when 16361 => pixel <= "000000";
      when 16362 => pixel <= "000000";
      when 16363 => pixel <= "000000";
      when 16364 => pixel <= "000000";
      when 16365 => pixel <= "000000";
      when 16366 => pixel <= "000000";
      when 16367 => pixel <= "000000";
      when 16368 => pixel <= "000000";
      when 16369 => pixel <= "000000";
      when 16370 => pixel <= "000000";
      when 16371 => pixel <= "000000";
      when 16372 => pixel <= "000000";
      when 16373 => pixel <= "000000";
      when 16374 => pixel <= "000000";
      when 16375 => pixel <= "000000";
      when 16376 => pixel <= "000000";
      when 16377 => pixel <= "000000";
      when 16378 => pixel <= "000000";
      when 16379 => pixel <= "000000";
      when 16380 => pixel <= "000000";
      when 16381 => pixel <= "000000";
      when 16382 => pixel <= "000000";
      when 16383 => pixel <= "000000";
      when 16384 => pixel <= "000000";
      when 16385 => pixel <= "000000";
      when 16386 => pixel <= "000000";
      when 16387 => pixel <= "000000";
      when 16388 => pixel <= "000000";
      when 16389 => pixel <= "000000";
      when 16390 => pixel <= "000000";
      when 16391 => pixel <= "000000";
      when 16392 => pixel <= "000000";
      when 16393 => pixel <= "000000";
      when 16394 => pixel <= "000000";
      when 16395 => pixel <= "000000";
      when 16396 => pixel <= "000000";
      when 16397 => pixel <= "000000";
      when 16398 => pixel <= "000000";
      when 16399 => pixel <= "000000";
      when 16400 => pixel <= "000000";
      when 16401 => pixel <= "000000";
      when 16402 => pixel <= "000000";
      when 16403 => pixel <= "000000";
      when 16404 => pixel <= "000000";
      when 16405 => pixel <= "000000";
      when 16406 => pixel <= "000000";
      when 16407 => pixel <= "000000";
      when 16408 => pixel <= "000000";
      when 16409 => pixel <= "000000";
      when 16410 => pixel <= "000000";
      when 16411 => pixel <= "000000";
      when 16412 => pixel <= "000000";
      when 16413 => pixel <= "000000";
      when 16414 => pixel <= "000000";
      when 16415 => pixel <= "000000";
      when 16416 => pixel <= "000000";
      when 16417 => pixel <= "000000";
      when 16418 => pixel <= "000000";
      when 16419 => pixel <= "000000";
      when 16420 => pixel <= "000000";
      when 16421 => pixel <= "000000";
      when 16422 => pixel <= "000000";
      when 16423 => pixel <= "000000";
      when 16424 => pixel <= "000000";
      when 16425 => pixel <= "000000";
      when 16426 => pixel <= "000000";
      when 16427 => pixel <= "000000";
      when 16428 => pixel <= "000000";
      when 16429 => pixel <= "000000";
      when 16430 => pixel <= "000000";
      when 16431 => pixel <= "000000";
      when 16432 => pixel <= "000000";
      when 16433 => pixel <= "000000";
      when 16434 => pixel <= "000000";
      when 16435 => pixel <= "000000";
      when 16436 => pixel <= "000000";
      when 16437 => pixel <= "000000";
      when 16438 => pixel <= "000000";
      when 16439 => pixel <= "000000";
      when 16440 => pixel <= "000000";
      when 16441 => pixel <= "000000";
      when 16442 => pixel <= "000000";
      when 16443 => pixel <= "000000";
      when 16444 => pixel <= "000000";
      when 16445 => pixel <= "000000";
      when 16446 => pixel <= "000000";
      when 16447 => pixel <= "000000";
      when 16448 => pixel <= "000000";
      when 16449 => pixel <= "000000";
      when 16450 => pixel <= "000000";
      when 16451 => pixel <= "000000";
      when 16452 => pixel <= "000000";
      when 16453 => pixel <= "000000";
      when 16454 => pixel <= "000000";
      when 16455 => pixel <= "000000";
      when 16456 => pixel <= "000000";
      when 16457 => pixel <= "000000";
      when 16458 => pixel <= "000000";
      when 16459 => pixel <= "000000";
      when 16460 => pixel <= "000000";
      when 16461 => pixel <= "000000";
      when 16462 => pixel <= "000000";
      when 16463 => pixel <= "000000";
      when 16464 => pixel <= "000000";
      when 16465 => pixel <= "000000";
      when 16466 => pixel <= "000000";
      when 16467 => pixel <= "000000";
      when 16468 => pixel <= "000000";
      when 16469 => pixel <= "000000";
      when 16470 => pixel <= "000000";
      when 16471 => pixel <= "000000";
      when 16472 => pixel <= "000000";
      when 16473 => pixel <= "000000";
      when 16474 => pixel <= "000000";
      when 16475 => pixel <= "000000";
      when 16476 => pixel <= "000000";
      when 16477 => pixel <= "000000";
      when 16478 => pixel <= "000000";
      when 16479 => pixel <= "000000";
      when 16480 => pixel <= "000000";
      when 16481 => pixel <= "000000";
      when 16482 => pixel <= "000000";
      when 16483 => pixel <= "000000";
      when 16484 => pixel <= "000000";
      when 16485 => pixel <= "000000";
      when 16486 => pixel <= "000000";
      when 16487 => pixel <= "000000";
      when 16488 => pixel <= "000000";
      when 16489 => pixel <= "000000";
      when 16490 => pixel <= "000000";
      when 16491 => pixel <= "000000";
      when 16492 => pixel <= "000000";
      when 16493 => pixel <= "000000";
      when 16494 => pixel <= "000000";
      when 16495 => pixel <= "000000";
      when 16496 => pixel <= "000000";
      when 16497 => pixel <= "000000";
      when 16498 => pixel <= "000000";
      when 16499 => pixel <= "000000";
      when 16500 => pixel <= "000000";
      when 16501 => pixel <= "000000";
      when 16502 => pixel <= "000000";
      when 16503 => pixel <= "000000";
      when 16504 => pixel <= "000000";
      when 16505 => pixel <= "000000";
      when 16506 => pixel <= "000000";
      when 16507 => pixel <= "000000";
      when 16508 => pixel <= "000000";
      when 16509 => pixel <= "000000";
      when 16510 => pixel <= "000000";
      when 16511 => pixel <= "000000";
      when 16512 => pixel <= "000000";
      when 16513 => pixel <= "000000";
      when 16514 => pixel <= "000000";
      when 16515 => pixel <= "000000";
      when 16516 => pixel <= "000000";
      when 16517 => pixel <= "000000";
      when 16518 => pixel <= "000000";
      when 16519 => pixel <= "000000";
      when 16520 => pixel <= "000000";
      when 16521 => pixel <= "000000";
      when 16522 => pixel <= "000000";
      when 16523 => pixel <= "000000";
      when 16524 => pixel <= "000000";
      when 16525 => pixel <= "000000";
      when 16526 => pixel <= "000000";
      when 16527 => pixel <= "000000";
      when 16528 => pixel <= "000000";
      when 16529 => pixel <= "000000";
      when 16530 => pixel <= "000000";
      when 16531 => pixel <= "000000";
      when 16532 => pixel <= "000000";
      when 16533 => pixel <= "000000";
      when 16534 => pixel <= "000000";
      when 16535 => pixel <= "000000";
      when 16536 => pixel <= "000000";
      when 16537 => pixel <= "000000";
      when 16538 => pixel <= "000000";
      when 16539 => pixel <= "000000";
      when 16540 => pixel <= "000000";
      when 16541 => pixel <= "000000";
      when 16542 => pixel <= "000000";
      when 16543 => pixel <= "000000";
      when 16544 => pixel <= "000000";
      when 16545 => pixel <= "000000";
      when 16546 => pixel <= "000000";
      when 16547 => pixel <= "000000";
      when 16548 => pixel <= "000000";
      when 16549 => pixel <= "000000";
      when 16550 => pixel <= "000000";
      when 16551 => pixel <= "000000";
      when 16552 => pixel <= "000000";
      when 16553 => pixel <= "000000";
      when 16554 => pixel <= "000000";
      when 16555 => pixel <= "000000";
      when 16556 => pixel <= "000000";
      when 16557 => pixel <= "000000";
      when 16558 => pixel <= "000000";
      when 16559 => pixel <= "000000";
      when 16560 => pixel <= "000000";
      when 16561 => pixel <= "000000";
      when 16562 => pixel <= "000000";
      when 16563 => pixel <= "000000";
      when 16564 => pixel <= "000000";
      when 16565 => pixel <= "000000";
      when 16566 => pixel <= "000000";
      when 16567 => pixel <= "000000";
      when 16568 => pixel <= "000000";
      when 16569 => pixel <= "000000";
      when 16570 => pixel <= "000000";
      when 16571 => pixel <= "000000";
      when 16572 => pixel <= "000000";
      when 16573 => pixel <= "000000";
      when 16574 => pixel <= "000000";
      when 16575 => pixel <= "000000";
      when 16576 => pixel <= "000000";
      when 16577 => pixel <= "000000";
      when 16578 => pixel <= "000000";
      when 16579 => pixel <= "000000";
      when 16580 => pixel <= "000000";
      when 16581 => pixel <= "000000";
      when 16582 => pixel <= "000000";
      when 16583 => pixel <= "000000";
      when 16584 => pixel <= "000000";
      when 16585 => pixel <= "000000";
      when 16586 => pixel <= "000000";
      when 16587 => pixel <= "000000";
      when 16588 => pixel <= "000000";
      when 16589 => pixel <= "000000";
      when 16590 => pixel <= "000000";
      when 16591 => pixel <= "000000";
      when 16592 => pixel <= "000000";
      when 16593 => pixel <= "000000";
      when 16594 => pixel <= "000000";
      when 16595 => pixel <= "000000";
      when 16596 => pixel <= "000000";
      when 16597 => pixel <= "000000";
      when 16598 => pixel <= "000000";
      when 16599 => pixel <= "000000";
      when 16600 => pixel <= "000000";
      when 16601 => pixel <= "000000";
      when 16602 => pixel <= "000000";
      when 16603 => pixel <= "000000";
      when 16604 => pixel <= "000000";
      when 16605 => pixel <= "000000";
      when 16606 => pixel <= "000000";
      when 16607 => pixel <= "000000";
      when 16608 => pixel <= "000000";
      when 16609 => pixel <= "000000";
      when 16610 => pixel <= "000000";
      when 16611 => pixel <= "000000";
      when 16612 => pixel <= "000000";
      when 16613 => pixel <= "000000";
      when 16614 => pixel <= "000000";
      when 16615 => pixel <= "000000";
      when 16616 => pixel <= "000000";
      when 16617 => pixel <= "000000";
      when 16618 => pixel <= "000000";
      when 16619 => pixel <= "000000";
      when 16620 => pixel <= "000000";
      when 16621 => pixel <= "000000";
      when 16622 => pixel <= "000000";
      when 16623 => pixel <= "000000";
      when 16624 => pixel <= "000000";
      when 16625 => pixel <= "000000";
      when 16626 => pixel <= "000000";
      when 16627 => pixel <= "000000";
      when 16628 => pixel <= "000000";
      when 16629 => pixel <= "000000";
      when 16630 => pixel <= "000000";
      when 16631 => pixel <= "000000";
      when 16632 => pixel <= "000000";
      when 16633 => pixel <= "000000";
      when 16634 => pixel <= "000000";
      when 16635 => pixel <= "000000";
      when 16636 => pixel <= "000000";
      when 16637 => pixel <= "000000";
      when 16638 => pixel <= "000000";
      when 16639 => pixel <= "000000";
      when 16640 => pixel <= "000000";
      when 16641 => pixel <= "000000";
      when 16642 => pixel <= "000000";
      when 16643 => pixel <= "000000";
      when 16644 => pixel <= "000000";
      when 16645 => pixel <= "000000";
      when 16646 => pixel <= "000000";
      when 16647 => pixel <= "000000";
      when 16648 => pixel <= "000000";
      when 16649 => pixel <= "000000";
      when 16650 => pixel <= "000000";
      when 16651 => pixel <= "000000";
      when 16652 => pixel <= "000000";
      when 16653 => pixel <= "000000";
      when 16654 => pixel <= "000000";
      when 16655 => pixel <= "000000";
      when 16656 => pixel <= "000000";
      when 16657 => pixel <= "000000";
      when 16658 => pixel <= "000000";
      when 16659 => pixel <= "000000";
      when 16660 => pixel <= "000000";
      when 16661 => pixel <= "000000";
      when 16662 => pixel <= "000000";
      when 16663 => pixel <= "000000";
      when 16664 => pixel <= "000000";
      when 16665 => pixel <= "000000";
      when 16666 => pixel <= "000000";
      when 16667 => pixel <= "000000";
      when 16668 => pixel <= "000000";
      when 16669 => pixel <= "000000";
      when 16670 => pixel <= "000000";
      when 16671 => pixel <= "000000";
      when 16672 => pixel <= "000000";
      when 16673 => pixel <= "000000";
      when 16674 => pixel <= "000000";
      when 16675 => pixel <= "000000";
      when 16676 => pixel <= "000000";
      when 16677 => pixel <= "000000";
      when 16678 => pixel <= "000000";
      when 16679 => pixel <= "000000";
      when 16680 => pixel <= "000000";
      when 16681 => pixel <= "000000";
      when 16682 => pixel <= "000000";
      when 16683 => pixel <= "000000";
      when 16684 => pixel <= "000000";
      when 16685 => pixel <= "000000";
      when 16686 => pixel <= "000000";
      when 16687 => pixel <= "000000";
      when 16688 => pixel <= "000000";
      when 16689 => pixel <= "000000";
      when 16690 => pixel <= "000000";
      when 16691 => pixel <= "000000";
      when 16692 => pixel <= "000000";
      when 16693 => pixel <= "000000";
      when 16694 => pixel <= "000000";
      when 16695 => pixel <= "000000";
      when 16696 => pixel <= "000000";
      when 16697 => pixel <= "000000";
      when 16698 => pixel <= "000000";
      when 16699 => pixel <= "000000";
      when 16700 => pixel <= "000000";
      when 16701 => pixel <= "000000";
      when 16702 => pixel <= "000000";
      when 16703 => pixel <= "000000";
      when 16704 => pixel <= "000000";
      when 16705 => pixel <= "000000";
      when 16706 => pixel <= "000000";
      when 16707 => pixel <= "000000";
      when 16708 => pixel <= "000000";
      when 16709 => pixel <= "000000";
      when 16710 => pixel <= "000000";
      when 16711 => pixel <= "000000";
      when 16712 => pixel <= "000000";
      when 16713 => pixel <= "000000";
      when 16714 => pixel <= "000000";
      when 16715 => pixel <= "000000";
      when 16716 => pixel <= "000000";
      when 16717 => pixel <= "000000";
      when 16718 => pixel <= "000000";
      when 16719 => pixel <= "000000";
      when 16720 => pixel <= "000000";
      when 16721 => pixel <= "000000";
      when 16722 => pixel <= "000000";
      when 16723 => pixel <= "000000";
      when 16724 => pixel <= "000000";
      when 16725 => pixel <= "000000";
      when 16726 => pixel <= "000000";
      when 16727 => pixel <= "000000";
      when 16728 => pixel <= "000000";
      when 16729 => pixel <= "000000";
      when 16730 => pixel <= "000000";
      when 16731 => pixel <= "000000";
      when 16732 => pixel <= "000000";
      when 16733 => pixel <= "000000";
      when 16734 => pixel <= "000000";
      when 16735 => pixel <= "000000";
      when 16736 => pixel <= "000000";
      when 16737 => pixel <= "000000";
      when 16738 => pixel <= "000000";
      when 16739 => pixel <= "000000";
      when 16740 => pixel <= "000000";
      when 16741 => pixel <= "000000";
      when 16742 => pixel <= "000000";
      when 16743 => pixel <= "000000";
      when 16744 => pixel <= "000000";
      when 16745 => pixel <= "000000";
      when 16746 => pixel <= "000000";
      when 16747 => pixel <= "000000";
      when 16748 => pixel <= "000000";
      when 16749 => pixel <= "000000";
      when 16750 => pixel <= "000000";
      when 16751 => pixel <= "000000";
      when 16752 => pixel <= "000000";
      when 16753 => pixel <= "000000";
      when 16754 => pixel <= "000000";
      when 16755 => pixel <= "000000";
      when 16756 => pixel <= "000000";
      when 16757 => pixel <= "000000";
      when 16758 => pixel <= "000000";
      when 16759 => pixel <= "000000";
      when 16760 => pixel <= "000000";
      when 16761 => pixel <= "000000";
      when 16762 => pixel <= "000000";
      when 16763 => pixel <= "000000";
      when 16764 => pixel <= "000000";
      when 16765 => pixel <= "000000";
      when 16766 => pixel <= "000000";
      when 16767 => pixel <= "000000";
      when 16768 => pixel <= "000000";
      when 16769 => pixel <= "000000";
      when 16770 => pixel <= "000000";
      when 16771 => pixel <= "000000";
      when 16772 => pixel <= "000000";
      when 16773 => pixel <= "000000";
      when 16774 => pixel <= "000000";
      when 16775 => pixel <= "000000";
      when 16776 => pixel <= "000000";
      when 16777 => pixel <= "000000";
      when 16778 => pixel <= "000000";
      when 16779 => pixel <= "000000";
      when 16780 => pixel <= "000000";
      when 16781 => pixel <= "000000";
      when 16782 => pixel <= "000000";
      when 16783 => pixel <= "000000";
      when 16784 => pixel <= "000000";
      when 16785 => pixel <= "000000";
      when 16786 => pixel <= "000000";
      when 16787 => pixel <= "000000";
      when 16788 => pixel <= "000000";
      when 16789 => pixel <= "000000";
      when 16790 => pixel <= "000000";
      when 16791 => pixel <= "000000";
      when 16792 => pixel <= "000000";
      when 16793 => pixel <= "000000";
      when 16794 => pixel <= "000000";
      when 16795 => pixel <= "000000";
      when 16796 => pixel <= "000000";
      when 16797 => pixel <= "000000";
      when 16798 => pixel <= "000000";
      when 16799 => pixel <= "000000";
      when 16800 => pixel <= "000000";
      when 16801 => pixel <= "000000";
      when 16802 => pixel <= "000000";
      when 16803 => pixel <= "000000";
      when 16804 => pixel <= "000000";
      when 16805 => pixel <= "000000";
      when 16806 => pixel <= "000000";
      when 16807 => pixel <= "000000";
      when 16808 => pixel <= "000000";
      when 16809 => pixel <= "000000";
      when 16810 => pixel <= "000000";
      when 16811 => pixel <= "000000";
      when 16812 => pixel <= "000000";
      when 16813 => pixel <= "000000";
      when 16814 => pixel <= "000000";
      when 16815 => pixel <= "000000";
      when 16816 => pixel <= "000000";
      when 16817 => pixel <= "000000";
      when 16818 => pixel <= "000000";
      when 16819 => pixel <= "000000";
      when 16820 => pixel <= "000000";
      when 16821 => pixel <= "000000";
      when 16822 => pixel <= "000000";
      when 16823 => pixel <= "000000";
      when 16824 => pixel <= "000000";
      when 16825 => pixel <= "000000";
      when 16826 => pixel <= "000000";
      when 16827 => pixel <= "000000";
      when 16828 => pixel <= "000000";
      when 16829 => pixel <= "000000";
      when 16830 => pixel <= "000000";
      when 16831 => pixel <= "000000";
      when 16832 => pixel <= "000000";
      when 16833 => pixel <= "000000";
      when 16834 => pixel <= "000000";
      when 16835 => pixel <= "000000";
      when 16836 => pixel <= "000000";
      when 16837 => pixel <= "000000";
      when 16838 => pixel <= "000000";
      when 16839 => pixel <= "000000";
      when 16840 => pixel <= "000000";
      when 16841 => pixel <= "000000";
      when 16842 => pixel <= "000000";
      when 16843 => pixel <= "000000";
      when 16844 => pixel <= "000000";
      when 16845 => pixel <= "000000";
      when 16846 => pixel <= "000000";
      when 16847 => pixel <= "000000";
      when 16848 => pixel <= "000000";
      when 16849 => pixel <= "000000";
      when 16850 => pixel <= "000000";
      when 16851 => pixel <= "000000";
      when 16852 => pixel <= "000000";
      when 16853 => pixel <= "000000";
      when 16854 => pixel <= "000000";
      when 16855 => pixel <= "000000";
      when 16856 => pixel <= "000000";
      when 16857 => pixel <= "000000";
      when 16858 => pixel <= "000000";
      when 16859 => pixel <= "000000";
      when 16860 => pixel <= "000000";
      when 16861 => pixel <= "000000";
      when 16862 => pixel <= "000000";
      when 16863 => pixel <= "000000";
      when 16864 => pixel <= "000000";
      when 16865 => pixel <= "000000";
      when 16866 => pixel <= "000000";
      when 16867 => pixel <= "000000";
      when 16868 => pixel <= "000000";
      when 16869 => pixel <= "000000";
      when 16870 => pixel <= "000000";
      when 16871 => pixel <= "000000";
      when 16872 => pixel <= "000000";
      when 16873 => pixel <= "000000";
      when 16874 => pixel <= "000000";
      when 16875 => pixel <= "000000";
      when 16876 => pixel <= "000000";
      when 16877 => pixel <= "000000";
      when 16878 => pixel <= "000000";
      when 16879 => pixel <= "000000";
      when 16880 => pixel <= "000000";
      when 16881 => pixel <= "000000";
      when 16882 => pixel <= "000000";
      when 16883 => pixel <= "000000";
      when 16884 => pixel <= "000000";
      when 16885 => pixel <= "000000";
      when 16886 => pixel <= "000000";
      when 16887 => pixel <= "000000";
      when 16888 => pixel <= "000000";
      when 16889 => pixel <= "000000";
      when 16890 => pixel <= "000000";
      when 16891 => pixel <= "000000";
      when 16892 => pixel <= "000000";
      when 16893 => pixel <= "000000";
      when 16894 => pixel <= "000000";
      when 16895 => pixel <= "000000";
      when 16896 => pixel <= "000000";
      when 16897 => pixel <= "000000";
      when 16898 => pixel <= "000000";
      when 16899 => pixel <= "000000";
      when 16900 => pixel <= "000000";
      when 16901 => pixel <= "000000";
      when 16902 => pixel <= "000000";
      when 16903 => pixel <= "000000";
      when 16904 => pixel <= "000000";
      when 16905 => pixel <= "000000";
      when 16906 => pixel <= "000000";
      when 16907 => pixel <= "000000";
      when 16908 => pixel <= "000000";
      when 16909 => pixel <= "000000";
      when 16910 => pixel <= "000000";
      when 16911 => pixel <= "000000";
      when 16912 => pixel <= "000000";
      when 16913 => pixel <= "000000";
      when 16914 => pixel <= "000000";
      when 16915 => pixel <= "000000";
      when 16916 => pixel <= "000000";
      when 16917 => pixel <= "000000";
      when 16918 => pixel <= "000000";
      when 16919 => pixel <= "000000";
      when 16920 => pixel <= "000000";
      when 16921 => pixel <= "000000";
      when 16922 => pixel <= "000000";
      when 16923 => pixel <= "000000";
      when 16924 => pixel <= "000000";
      when 16925 => pixel <= "000000";
      when 16926 => pixel <= "000000";
      when 16927 => pixel <= "000000";
      when 16928 => pixel <= "000000";
      when 16929 => pixel <= "000000";
      when 16930 => pixel <= "000000";
      when 16931 => pixel <= "000000";
      when 16932 => pixel <= "000000";
      when 16933 => pixel <= "000000";
      when 16934 => pixel <= "000000";
      when 16935 => pixel <= "000000";
      when 16936 => pixel <= "000000";
      when 16937 => pixel <= "000000";
      when 16938 => pixel <= "000000";
      when 16939 => pixel <= "000000";
      when 16940 => pixel <= "000000";
      when 16941 => pixel <= "000000";
      when 16942 => pixel <= "000000";
      when 16943 => pixel <= "000000";
      when 16944 => pixel <= "000000";
      when 16945 => pixel <= "000000";
      when 16946 => pixel <= "000000";
      when 16947 => pixel <= "000000";
      when 16948 => pixel <= "000000";
      when 16949 => pixel <= "000000";
      when 16950 => pixel <= "000000";
      when 16951 => pixel <= "000000";
      when 16952 => pixel <= "000000";
      when 16953 => pixel <= "000000";
      when 16954 => pixel <= "000000";
      when 16955 => pixel <= "000000";
      when 16956 => pixel <= "000000";
      when 16957 => pixel <= "000000";
      when 16958 => pixel <= "000000";
      when 16959 => pixel <= "000000";
      when 16960 => pixel <= "000000";
      when 16961 => pixel <= "000000";
      when 16962 => pixel <= "000000";
      when 16963 => pixel <= "000000";
      when 16964 => pixel <= "000000";
      when 16965 => pixel <= "000000";
      when 16966 => pixel <= "000000";
      when 16967 => pixel <= "000000";
      when 16968 => pixel <= "000000";
      when 16969 => pixel <= "000000";
      when 16970 => pixel <= "000000";
      when 16971 => pixel <= "000000";
      when 16972 => pixel <= "000000";
      when 16973 => pixel <= "000000";
      when 16974 => pixel <= "000000";
      when 16975 => pixel <= "000000";
      when 16976 => pixel <= "000000";
      when 16977 => pixel <= "000000";
      when 16978 => pixel <= "000000";
      when 16979 => pixel <= "000000";
      when 16980 => pixel <= "000000";
      when 16981 => pixel <= "000000";
      when 16982 => pixel <= "000000";
      when 16983 => pixel <= "000000";
      when 16984 => pixel <= "000000";
      when 16985 => pixel <= "000000";
      when 16986 => pixel <= "000000";
      when 16987 => pixel <= "000000";
      when 16988 => pixel <= "000000";
      when 16989 => pixel <= "000000";
      when 16990 => pixel <= "000000";
      when 16991 => pixel <= "000000";
      when 16992 => pixel <= "000000";
      when 16993 => pixel <= "000000";
      when 16994 => pixel <= "000000";
      when 16995 => pixel <= "000000";
      when 16996 => pixel <= "000000";
      when 16997 => pixel <= "000000";
      when 16998 => pixel <= "000000";
      when 16999 => pixel <= "000000";
      when 17000 => pixel <= "000000";
      when 17001 => pixel <= "000000";
      when 17002 => pixel <= "000000";
      when 17003 => pixel <= "000000";
      when 17004 => pixel <= "000000";
      when 17005 => pixel <= "000000";
      when 17006 => pixel <= "000000";
      when 17007 => pixel <= "000000";
      when 17008 => pixel <= "000000";
      when 17009 => pixel <= "000000";
      when 17010 => pixel <= "000000";
      when 17011 => pixel <= "000000";
      when 17012 => pixel <= "000000";
      when 17013 => pixel <= "000000";
      when 17014 => pixel <= "000000";
      when 17015 => pixel <= "000000";
      when 17016 => pixel <= "000000";
      when 17017 => pixel <= "000000";
      when 17018 => pixel <= "000000";
      when 17019 => pixel <= "000000";
      when 17020 => pixel <= "000000";
      when 17021 => pixel <= "000000";
      when 17022 => pixel <= "000000";
      when 17023 => pixel <= "000000";
      when 17024 => pixel <= "000000";
      when 17025 => pixel <= "000000";
      when 17026 => pixel <= "000000";
      when 17027 => pixel <= "000000";
      when 17028 => pixel <= "000000";
      when 17029 => pixel <= "000000";
      when 17030 => pixel <= "000000";
      when 17031 => pixel <= "000000";
      when 17032 => pixel <= "000000";
      when 17033 => pixel <= "000000";
      when 17034 => pixel <= "000000";
      when 17035 => pixel <= "000000";
      when 17036 => pixel <= "000000";
      when 17037 => pixel <= "000000";
      when 17038 => pixel <= "000000";
      when 17039 => pixel <= "000000";
      when 17040 => pixel <= "000000";
      when 17041 => pixel <= "000000";
      when 17042 => pixel <= "000000";
      when 17043 => pixel <= "000000";
      when 17044 => pixel <= "000000";
      when 17045 => pixel <= "000000";
      when 17046 => pixel <= "000000";
      when 17047 => pixel <= "000000";
      when 17048 => pixel <= "000000";
      when 17049 => pixel <= "000000";
      when 17050 => pixel <= "000000";
      when 17051 => pixel <= "000000";
      when 17052 => pixel <= "000000";
      when 17053 => pixel <= "000000";
      when 17054 => pixel <= "000000";
      when 17055 => pixel <= "000000";
      when 17056 => pixel <= "000000";
      when 17057 => pixel <= "000000";
      when 17058 => pixel <= "000000";
      when 17059 => pixel <= "000000";
      when 17060 => pixel <= "000000";
      when 17061 => pixel <= "000000";
      when 17062 => pixel <= "000000";
      when 17063 => pixel <= "000000";
      when 17064 => pixel <= "000000";
      when 17065 => pixel <= "000000";
      when 17066 => pixel <= "000000";
      when 17067 => pixel <= "000000";
      when 17068 => pixel <= "000000";
      when 17069 => pixel <= "000000";
      when 17070 => pixel <= "000000";
      when 17071 => pixel <= "000000";
      when 17072 => pixel <= "000000";
      when 17073 => pixel <= "000000";
      when 17074 => pixel <= "000000";
      when 17075 => pixel <= "000000";
      when 17076 => pixel <= "000000";
      when 17077 => pixel <= "000000";
      when 17078 => pixel <= "000000";
      when 17079 => pixel <= "000000";
      when 17080 => pixel <= "000000";
      when 17081 => pixel <= "000000";
      when 17082 => pixel <= "000000";
      when 17083 => pixel <= "000000";
      when 17084 => pixel <= "000000";
      when 17085 => pixel <= "000000";
      when 17086 => pixel <= "000000";
      when 17087 => pixel <= "000000";
      when 17088 => pixel <= "000000";
      when 17089 => pixel <= "000000";
      when 17090 => pixel <= "000000";
      when 17091 => pixel <= "000000";
      when 17092 => pixel <= "000000";
      when 17093 => pixel <= "000000";
      when 17094 => pixel <= "000000";
      when 17095 => pixel <= "000000";
      when 17096 => pixel <= "000000";
      when 17097 => pixel <= "000000";
      when 17098 => pixel <= "000000";
      when 17099 => pixel <= "000000";
      when 17100 => pixel <= "000000";
      when 17101 => pixel <= "000000";
      when 17102 => pixel <= "000000";
      when 17103 => pixel <= "000000";
      when 17104 => pixel <= "000000";
      when 17105 => pixel <= "000000";
      when 17106 => pixel <= "000000";
      when 17107 => pixel <= "000000";
      when 17108 => pixel <= "000000";
      when 17109 => pixel <= "000000";
      when 17110 => pixel <= "000000";
      when 17111 => pixel <= "000000";
      when 17112 => pixel <= "000000";
      when 17113 => pixel <= "000000";
      when 17114 => pixel <= "000000";
      when 17115 => pixel <= "000000";
      when 17116 => pixel <= "000000";
      when 17117 => pixel <= "000000";
      when 17118 => pixel <= "000000";
      when 17119 => pixel <= "000000";
      when 17120 => pixel <= "000000";
      when 17121 => pixel <= "000000";
      when 17122 => pixel <= "000000";
      when 17123 => pixel <= "000000";
      when 17124 => pixel <= "000000";
      when 17125 => pixel <= "000000";
      when 17126 => pixel <= "000000";
      when 17127 => pixel <= "000000";
      when 17128 => pixel <= "000000";
      when 17129 => pixel <= "000000";
      when 17130 => pixel <= "000000";
      when 17131 => pixel <= "000000";
      when 17132 => pixel <= "000000";
      when 17133 => pixel <= "000000";
      when 17134 => pixel <= "000000";
      when 17135 => pixel <= "000000";
      when 17136 => pixel <= "000000";
      when 17137 => pixel <= "000000";
      when 17138 => pixel <= "000000";
      when 17139 => pixel <= "000000";
      when 17140 => pixel <= "000000";
      when 17141 => pixel <= "000000";
      when 17142 => pixel <= "000000";
      when 17143 => pixel <= "000000";
      when 17144 => pixel <= "000000";
      when 17145 => pixel <= "000000";
      when 17146 => pixel <= "000000";
      when 17147 => pixel <= "000000";
      when 17148 => pixel <= "000000";
      when 17149 => pixel <= "000000";
      when 17150 => pixel <= "000000";
      when 17151 => pixel <= "000000";
      when 17152 => pixel <= "000000";
      when 17153 => pixel <= "000000";
      when 17154 => pixel <= "000000";
      when 17155 => pixel <= "000000";
      when 17156 => pixel <= "000000";
      when 17157 => pixel <= "000000";
      when 17158 => pixel <= "000000";
      when 17159 => pixel <= "000000";
      when 17160 => pixel <= "000000";
      when 17161 => pixel <= "000000";
      when 17162 => pixel <= "000000";
      when 17163 => pixel <= "000000";
      when 17164 => pixel <= "000000";
      when 17165 => pixel <= "000000";
      when 17166 => pixel <= "000000";
      when 17167 => pixel <= "000000";
      when 17168 => pixel <= "000000";
      when 17169 => pixel <= "000000";
      when 17170 => pixel <= "000000";
      when 17171 => pixel <= "000000";
      when 17172 => pixel <= "000000";
      when 17173 => pixel <= "000000";
      when 17174 => pixel <= "000000";
      when 17175 => pixel <= "000000";
      when 17176 => pixel <= "000000";
      when 17177 => pixel <= "000000";
      when 17178 => pixel <= "000000";
      when 17179 => pixel <= "000000";
      when 17180 => pixel <= "000000";
      when 17181 => pixel <= "000000";
      when 17182 => pixel <= "000000";
      when 17183 => pixel <= "000000";
      when 17184 => pixel <= "000000";
      when 17185 => pixel <= "000000";
      when 17186 => pixel <= "000000";
      when 17187 => pixel <= "000000";
      when 17188 => pixel <= "000000";
      when 17189 => pixel <= "000000";
      when 17190 => pixel <= "000000";
      when 17191 => pixel <= "000000";
      when 17192 => pixel <= "000000";
      when 17193 => pixel <= "000000";
      when 17194 => pixel <= "000000";
      when 17195 => pixel <= "000000";
      when 17196 => pixel <= "000000";
      when 17197 => pixel <= "000000";
      when 17198 => pixel <= "000000";
      when 17199 => pixel <= "000000";
      when 17200 => pixel <= "000000";
      when 17201 => pixel <= "000000";
      when 17202 => pixel <= "000000";
      when 17203 => pixel <= "000000";
      when 17204 => pixel <= "000000";
      when 17205 => pixel <= "000000";
      when 17206 => pixel <= "000000";
      when 17207 => pixel <= "000000";
      when 17208 => pixel <= "000000";
      when 17209 => pixel <= "000000";
      when 17210 => pixel <= "000000";
      when 17211 => pixel <= "000000";
      when 17212 => pixel <= "000000";
      when 17213 => pixel <= "000000";
      when 17214 => pixel <= "000000";
      when 17215 => pixel <= "000000";
      when 17216 => pixel <= "000000";
      when 17217 => pixel <= "000000";
      when 17218 => pixel <= "000000";
      when 17219 => pixel <= "000000";
      when 17220 => pixel <= "000000";
      when 17221 => pixel <= "000000";
      when 17222 => pixel <= "000000";
      when 17223 => pixel <= "000000";
      when 17224 => pixel <= "000000";
      when 17225 => pixel <= "000000";
      when 17226 => pixel <= "000000";
      when 17227 => pixel <= "000000";
      when 17228 => pixel <= "000000";
      when 17229 => pixel <= "000000";
      when 17230 => pixel <= "000000";
      when 17231 => pixel <= "000000";
      when 17232 => pixel <= "000000";
      when 17233 => pixel <= "000000";
      when 17234 => pixel <= "000000";
      when 17235 => pixel <= "000000";
      when 17236 => pixel <= "000000";
      when 17237 => pixel <= "000000";
      when 17238 => pixel <= "000000";
      when 17239 => pixel <= "000000";
      when 17240 => pixel <= "000000";
      when 17241 => pixel <= "000000";
      when 17242 => pixel <= "000000";
      when 17243 => pixel <= "000000";
      when 17244 => pixel <= "000000";
      when 17245 => pixel <= "000000";
      when 17246 => pixel <= "000000";
      when 17247 => pixel <= "000000";
      when 17248 => pixel <= "000000";
      when 17249 => pixel <= "000000";
      when 17250 => pixel <= "000000";
      when 17251 => pixel <= "000000";
      when 17252 => pixel <= "000000";
      when 17253 => pixel <= "000000";
      when 17254 => pixel <= "000000";
      when 17255 => pixel <= "000000";
      when 17256 => pixel <= "000000";
      when 17257 => pixel <= "000000";
      when 17258 => pixel <= "000000";
      when 17259 => pixel <= "000000";
      when 17260 => pixel <= "000000";
      when 17261 => pixel <= "000000";
      when 17262 => pixel <= "000000";
      when 17263 => pixel <= "000000";
      when 17264 => pixel <= "000000";
      when 17265 => pixel <= "000000";
      when 17266 => pixel <= "000000";
      when 17267 => pixel <= "000000";
      when 17268 => pixel <= "000000";
      when 17269 => pixel <= "000000";
      when 17270 => pixel <= "000000";
      when 17271 => pixel <= "000000";
      when 17272 => pixel <= "000000";
      when 17273 => pixel <= "000000";
      when 17274 => pixel <= "000000";
      when 17275 => pixel <= "000000";
      when 17276 => pixel <= "000000";
      when 17277 => pixel <= "000000";
      when 17278 => pixel <= "000000";
      when 17279 => pixel <= "000000";
      when 17280 => pixel <= "000000";
      when 17281 => pixel <= "000000";
      when 17282 => pixel <= "000000";
      when 17283 => pixel <= "000000";
      when 17284 => pixel <= "000000";
      when 17285 => pixel <= "000000";
      when 17286 => pixel <= "000000";
      when 17287 => pixel <= "000000";
      when 17288 => pixel <= "000000";
      when 17289 => pixel <= "000000";
      when 17290 => pixel <= "000000";
      when 17291 => pixel <= "000000";
      when 17292 => pixel <= "000000";
      when 17293 => pixel <= "000000";
      when 17294 => pixel <= "000000";
      when 17295 => pixel <= "000000";
      when 17296 => pixel <= "000000";
      when 17297 => pixel <= "000000";
      when 17298 => pixel <= "000000";
      when 17299 => pixel <= "000000";
      when 17300 => pixel <= "000000";
      when 17301 => pixel <= "000000";
      when 17302 => pixel <= "000000";
      when 17303 => pixel <= "000000";
      when 17304 => pixel <= "000000";
      when 17305 => pixel <= "000000";
      when 17306 => pixel <= "000000";
      when 17307 => pixel <= "000000";
      when 17308 => pixel <= "000000";
      when 17309 => pixel <= "000000";
      when 17310 => pixel <= "000000";
      when 17311 => pixel <= "000000";
      when 17312 => pixel <= "000000";
      when 17313 => pixel <= "000000";
      when 17314 => pixel <= "000000";
      when 17315 => pixel <= "000000";
      when 17316 => pixel <= "000000";
      when 17317 => pixel <= "000000";
      when 17318 => pixel <= "000000";
      when 17319 => pixel <= "000000";
      when 17320 => pixel <= "000000";
      when 17321 => pixel <= "000000";
      when 17322 => pixel <= "000000";
      when 17323 => pixel <= "000000";
      when 17324 => pixel <= "000000";
      when 17325 => pixel <= "000000";
      when 17326 => pixel <= "000000";
      when 17327 => pixel <= "000000";
      when 17328 => pixel <= "000000";
      when 17329 => pixel <= "000000";
      when 17330 => pixel <= "000000";
      when 17331 => pixel <= "000000";
      when 17332 => pixel <= "000000";
      when 17333 => pixel <= "000000";
      when 17334 => pixel <= "000000";
      when 17335 => pixel <= "000000";
      when 17336 => pixel <= "000000";
      when 17337 => pixel <= "000000";
      when 17338 => pixel <= "000000";
      when 17339 => pixel <= "000000";
      when 17340 => pixel <= "000000";
      when 17341 => pixel <= "000000";
      when 17342 => pixel <= "000000";
      when 17343 => pixel <= "000000";
      when 17344 => pixel <= "000000";
      when 17345 => pixel <= "000000";
      when 17346 => pixel <= "000000";
      when 17347 => pixel <= "000000";
      when 17348 => pixel <= "000000";
      when 17349 => pixel <= "000000";
      when 17350 => pixel <= "000000";
      when 17351 => pixel <= "000000";
      when 17352 => pixel <= "000000";
      when 17353 => pixel <= "000000";
      when 17354 => pixel <= "000000";
      when 17355 => pixel <= "000000";
      when 17356 => pixel <= "000000";
      when 17357 => pixel <= "000000";
      when 17358 => pixel <= "000000";
      when 17359 => pixel <= "000000";
      when 17360 => pixel <= "000000";
      when 17361 => pixel <= "000000";
      when 17362 => pixel <= "000000";
      when 17363 => pixel <= "000000";
      when 17364 => pixel <= "000000";
      when 17365 => pixel <= "000000";
      when 17366 => pixel <= "000000";
      when 17367 => pixel <= "000000";
      when 17368 => pixel <= "000000";
      when 17369 => pixel <= "000000";
      when 17370 => pixel <= "000000";
      when 17371 => pixel <= "000000";
      when 17372 => pixel <= "000000";
      when 17373 => pixel <= "000000";
      when 17374 => pixel <= "000000";
      when 17375 => pixel <= "000000";
      when 17376 => pixel <= "000000";
      when 17377 => pixel <= "000000";
      when 17378 => pixel <= "000000";
      when 17379 => pixel <= "000000";
      when 17380 => pixel <= "000000";
      when 17381 => pixel <= "000000";
      when 17382 => pixel <= "000000";
      when 17383 => pixel <= "000000";
      when 17384 => pixel <= "000000";
      when 17385 => pixel <= "000000";
      when 17386 => pixel <= "000000";
      when 17387 => pixel <= "000000";
      when 17388 => pixel <= "000000";
      when 17389 => pixel <= "000000";
      when 17390 => pixel <= "000000";
      when 17391 => pixel <= "000000";
      when 17392 => pixel <= "000000";
      when 17393 => pixel <= "000000";
      when 17394 => pixel <= "000000";
      when 17395 => pixel <= "000000";
      when 17396 => pixel <= "000000";
      when 17397 => pixel <= "000000";
      when 17398 => pixel <= "000000";
      when 17399 => pixel <= "000000";
      when 17400 => pixel <= "000000";
      when 17401 => pixel <= "000000";
      when 17402 => pixel <= "000000";
      when 17403 => pixel <= "000000";
      when 17404 => pixel <= "000000";
      when 17405 => pixel <= "000000";
      when 17406 => pixel <= "000000";
      when 17407 => pixel <= "000000";
      when 17408 => pixel <= "000000";
      when 17409 => pixel <= "000000";
      when 17410 => pixel <= "000000";
      when 17411 => pixel <= "000000";
      when 17412 => pixel <= "000000";
      when 17413 => pixel <= "000000";
      when 17414 => pixel <= "000000";
      when 17415 => pixel <= "000000";
      when 17416 => pixel <= "000000";
      when 17417 => pixel <= "000000";
      when 17418 => pixel <= "000000";
      when 17419 => pixel <= "000000";
      when 17420 => pixel <= "000000";
      when 17421 => pixel <= "000000";
      when 17422 => pixel <= "000000";
      when 17423 => pixel <= "000000";
      when 17424 => pixel <= "000000";
      when 17425 => pixel <= "000000";
      when 17426 => pixel <= "000000";
      when 17427 => pixel <= "000000";
      when 17428 => pixel <= "000000";
      when 17429 => pixel <= "000000";
      when 17430 => pixel <= "000000";
      when 17431 => pixel <= "000000";
      when 17432 => pixel <= "000000";
      when 17433 => pixel <= "000000";
      when 17434 => pixel <= "000000";
      when 17435 => pixel <= "000000";
      when 17436 => pixel <= "000000";
      when 17437 => pixel <= "000000";
      when 17438 => pixel <= "000000";
      when 17439 => pixel <= "000000";
      when 17440 => pixel <= "000000";
      when 17441 => pixel <= "000000";
      when 17442 => pixel <= "000000";
      when 17443 => pixel <= "000000";
      when 17444 => pixel <= "000000";
      when 17445 => pixel <= "000000";
      when 17446 => pixel <= "000000";
      when 17447 => pixel <= "000000";
      when 17448 => pixel <= "000000";
      when 17449 => pixel <= "000000";
      when 17450 => pixel <= "000000";
      when 17451 => pixel <= "000000";
      when 17452 => pixel <= "000000";
      when 17453 => pixel <= "000000";
      when 17454 => pixel <= "000000";
      when 17455 => pixel <= "000000";
      when 17456 => pixel <= "000000";
      when 17457 => pixel <= "000000";
      when 17458 => pixel <= "000000";
      when 17459 => pixel <= "000000";
      when 17460 => pixel <= "000000";
      when 17461 => pixel <= "000000";
      when 17462 => pixel <= "000000";
      when 17463 => pixel <= "000000";
      when 17464 => pixel <= "000000";
      when 17465 => pixel <= "000000";
      when 17466 => pixel <= "000000";
      when 17467 => pixel <= "000000";
      when 17468 => pixel <= "000000";
      when 17469 => pixel <= "000000";
      when 17470 => pixel <= "000000";
      when 17471 => pixel <= "000000";
      when 17472 => pixel <= "000000";
      when 17473 => pixel <= "000000";
      when 17474 => pixel <= "000000";
      when 17475 => pixel <= "000000";
      when 17476 => pixel <= "000000";
      when 17477 => pixel <= "000000";
      when 17478 => pixel <= "000000";
      when 17479 => pixel <= "000000";
      when 17480 => pixel <= "000000";
      when 17481 => pixel <= "000000";
      when 17482 => pixel <= "000000";
      when 17483 => pixel <= "000000";
      when 17484 => pixel <= "000000";
      when 17485 => pixel <= "000000";
      when 17486 => pixel <= "000000";
      when 17487 => pixel <= "000000";
      when 17488 => pixel <= "000000";
      when 17489 => pixel <= "000000";
      when 17490 => pixel <= "000000";
      when 17491 => pixel <= "000000";
      when 17492 => pixel <= "000000";
      when 17493 => pixel <= "000000";
      when 17494 => pixel <= "000000";
      when 17495 => pixel <= "000000";
      when 17496 => pixel <= "000000";
      when 17497 => pixel <= "000000";
      when 17498 => pixel <= "000000";
      when 17499 => pixel <= "000000";
      when 17500 => pixel <= "000000";
      when 17501 => pixel <= "000000";
      when 17502 => pixel <= "000000";
      when 17503 => pixel <= "000000";
      when 17504 => pixel <= "000000";
      when 17505 => pixel <= "000000";
      when 17506 => pixel <= "000000";
      when 17507 => pixel <= "000000";
      when 17508 => pixel <= "000000";
      when 17509 => pixel <= "000000";
      when 17510 => pixel <= "000000";
      when 17511 => pixel <= "000000";
      when 17512 => pixel <= "000000";
      when 17513 => pixel <= "000000";
      when 17514 => pixel <= "000000";
      when 17515 => pixel <= "000000";
      when 17516 => pixel <= "000000";
      when 17517 => pixel <= "000000";
      when 17518 => pixel <= "000000";
      when 17519 => pixel <= "000000";
      when 17520 => pixel <= "000000";
      when 17521 => pixel <= "000000";
      when 17522 => pixel <= "000000";
      when 17523 => pixel <= "000000";
      when 17524 => pixel <= "000000";
      when 17525 => pixel <= "000000";
      when 17526 => pixel <= "000000";
      when 17527 => pixel <= "000000";
      when 17528 => pixel <= "000000";
      when 17529 => pixel <= "000000";
      when 17530 => pixel <= "000000";
      when 17531 => pixel <= "000000";
      when 17532 => pixel <= "000000";
      when 17533 => pixel <= "000000";
      when 17534 => pixel <= "000000";
      when 17535 => pixel <= "000000";
      when 17536 => pixel <= "000000";
      when 17537 => pixel <= "000000";
      when 17538 => pixel <= "000000";
      when 17539 => pixel <= "000000";
      when 17540 => pixel <= "000000";
      when 17541 => pixel <= "000000";
      when 17542 => pixel <= "000000";
      when 17543 => pixel <= "000000";
      when 17544 => pixel <= "000000";
      when 17545 => pixel <= "000000";
      when 17546 => pixel <= "000000";
      when 17547 => pixel <= "000000";
      when 17548 => pixel <= "000000";
      when 17549 => pixel <= "000000";
      when 17550 => pixel <= "000000";
      when 17551 => pixel <= "000000";
      when 17552 => pixel <= "000000";
      when 17553 => pixel <= "000000";
      when 17554 => pixel <= "000000";
      when 17555 => pixel <= "000000";
      when 17556 => pixel <= "000000";
      when 17557 => pixel <= "000000";
      when 17558 => pixel <= "000000";
      when 17559 => pixel <= "000000";
      when 17560 => pixel <= "000000";
      when 17561 => pixel <= "000000";
      when 17562 => pixel <= "000000";
      when 17563 => pixel <= "000000";
      when 17564 => pixel <= "000000";
      when 17565 => pixel <= "000000";
      when 17566 => pixel <= "000000";
      when 17567 => pixel <= "000000";
      when 17568 => pixel <= "000000";
      when 17569 => pixel <= "000000";
      when 17570 => pixel <= "000000";
      when 17571 => pixel <= "000000";
      when 17572 => pixel <= "000000";
      when 17573 => pixel <= "000000";
      when 17574 => pixel <= "000000";
      when 17575 => pixel <= "000000";
      when 17576 => pixel <= "000000";
      when 17577 => pixel <= "000000";
      when 17578 => pixel <= "000000";
      when 17579 => pixel <= "000000";
      when 17580 => pixel <= "000000";
      when 17581 => pixel <= "000000";
      when 17582 => pixel <= "000000";
      when 17583 => pixel <= "000000";
      when 17584 => pixel <= "000000";
      when 17585 => pixel <= "000000";
      when 17586 => pixel <= "000000";
      when 17587 => pixel <= "000000";
      when 17588 => pixel <= "000000";
      when 17589 => pixel <= "000000";
      when 17590 => pixel <= "000000";
      when 17591 => pixel <= "000000";
      when 17592 => pixel <= "000000";
      when 17593 => pixel <= "000000";
      when 17594 => pixel <= "000000";
      when 17595 => pixel <= "000000";
      when 17596 => pixel <= "000000";
      when 17597 => pixel <= "000000";
      when 17598 => pixel <= "000000";
      when 17599 => pixel <= "000000";
      when 17600 => pixel <= "000000";
      when 17601 => pixel <= "000000";
      when 17602 => pixel <= "000000";
      when 17603 => pixel <= "000000";
      when 17604 => pixel <= "000000";
      when 17605 => pixel <= "000000";
      when 17606 => pixel <= "000000";
      when 17607 => pixel <= "000000";
      when 17608 => pixel <= "000000";
      when 17609 => pixel <= "000000";
      when 17610 => pixel <= "000000";
      when 17611 => pixel <= "000000";
      when 17612 => pixel <= "000000";
      when 17613 => pixel <= "000000";
      when 17614 => pixel <= "000000";
      when 17615 => pixel <= "000000";
      when 17616 => pixel <= "000000";
      when 17617 => pixel <= "000000";
      when 17618 => pixel <= "000000";
      when 17619 => pixel <= "000000";
      when 17620 => pixel <= "000000";
      when 17621 => pixel <= "000000";
      when 17622 => pixel <= "000000";
      when 17623 => pixel <= "000000";
      when 17624 => pixel <= "000000";
      when 17625 => pixel <= "000000";
      when 17626 => pixel <= "000000";
      when 17627 => pixel <= "000000";
      when 17628 => pixel <= "000000";
      when 17629 => pixel <= "000000";
      when 17630 => pixel <= "000000";
      when 17631 => pixel <= "000000";
      when 17632 => pixel <= "000000";
      when 17633 => pixel <= "000000";
      when 17634 => pixel <= "000000";
      when 17635 => pixel <= "000000";
      when 17636 => pixel <= "000000";
      when 17637 => pixel <= "000000";
      when 17638 => pixel <= "000000";
      when 17639 => pixel <= "000000";
      when 17640 => pixel <= "000000";
      when 17641 => pixel <= "000000";
      when 17642 => pixel <= "000000";
      when 17643 => pixel <= "000000";
      when 17644 => pixel <= "000000";
      when 17645 => pixel <= "000000";
      when 17646 => pixel <= "000000";
      when 17647 => pixel <= "000000";
      when 17648 => pixel <= "000000";
      when 17649 => pixel <= "000000";
      when 17650 => pixel <= "000000";
      when 17651 => pixel <= "000000";
      when 17652 => pixel <= "000000";
      when 17653 => pixel <= "000000";
      when 17654 => pixel <= "000000";
      when 17655 => pixel <= "000000";
      when 17656 => pixel <= "000000";
      when 17657 => pixel <= "000000";
      when 17658 => pixel <= "000000";
      when 17659 => pixel <= "000000";
      when 17660 => pixel <= "000000";
      when 17661 => pixel <= "000000";
      when 17662 => pixel <= "000000";
      when 17663 => pixel <= "000000";
      when 17664 => pixel <= "000000";
      when 17665 => pixel <= "000000";
      when 17666 => pixel <= "000000";
      when 17667 => pixel <= "000000";
      when 17668 => pixel <= "000000";
      when 17669 => pixel <= "000000";
      when 17670 => pixel <= "000000";
      when 17671 => pixel <= "000000";
      when 17672 => pixel <= "000000";
      when 17673 => pixel <= "000000";
      when 17674 => pixel <= "000000";
      when 17675 => pixel <= "000000";
      when 17676 => pixel <= "000000";
      when 17677 => pixel <= "000000";
      when 17678 => pixel <= "000000";
      when 17679 => pixel <= "000000";
      when 17680 => pixel <= "000000";
      when 17681 => pixel <= "000000";
      when 17682 => pixel <= "000000";
      when 17683 => pixel <= "000000";
      when 17684 => pixel <= "000000";
      when 17685 => pixel <= "000000";
      when 17686 => pixel <= "000000";
      when 17687 => pixel <= "000000";
      when 17688 => pixel <= "000000";
      when 17689 => pixel <= "000000";
      when 17690 => pixel <= "000000";
      when 17691 => pixel <= "000000";
      when 17692 => pixel <= "000000";
      when 17693 => pixel <= "000000";
      when 17694 => pixel <= "000000";
      when 17695 => pixel <= "000000";
      when 17696 => pixel <= "000000";
      when 17697 => pixel <= "000000";
      when 17698 => pixel <= "000000";
      when 17699 => pixel <= "000000";
      when 17700 => pixel <= "000000";
      when 17701 => pixel <= "000000";
      when 17702 => pixel <= "000000";
      when 17703 => pixel <= "000000";
      when 17704 => pixel <= "000000";
      when 17705 => pixel <= "000000";
      when 17706 => pixel <= "000000";
      when 17707 => pixel <= "000000";
      when 17708 => pixel <= "000000";
      when 17709 => pixel <= "000000";
      when 17710 => pixel <= "000000";
      when 17711 => pixel <= "000000";
      when 17712 => pixel <= "000000";
      when 17713 => pixel <= "000000";
      when 17714 => pixel <= "000000";
      when 17715 => pixel <= "000000";
      when 17716 => pixel <= "000000";
      when 17717 => pixel <= "000000";
      when 17718 => pixel <= "000000";
      when 17719 => pixel <= "000000";
      when 17720 => pixel <= "000000";
      when 17721 => pixel <= "000000";
      when 17722 => pixel <= "000000";
      when 17723 => pixel <= "000000";
      when 17724 => pixel <= "000000";
      when 17725 => pixel <= "000000";
      when 17726 => pixel <= "000000";
      when 17727 => pixel <= "000000";
      when 17728 => pixel <= "000000";
      when 17729 => pixel <= "000000";
      when 17730 => pixel <= "000000";
      when 17731 => pixel <= "000000";
      when 17732 => pixel <= "000000";
      when 17733 => pixel <= "000000";
      when 17734 => pixel <= "000000";
      when 17735 => pixel <= "000000";
      when 17736 => pixel <= "000000";
      when 17737 => pixel <= "000000";
      when 17738 => pixel <= "000000";
      when 17739 => pixel <= "000000";
      when 17740 => pixel <= "000000";
      when 17741 => pixel <= "000000";
      when 17742 => pixel <= "000000";
      when 17743 => pixel <= "000000";
      when 17744 => pixel <= "000000";
      when 17745 => pixel <= "000000";
      when 17746 => pixel <= "000000";
      when 17747 => pixel <= "000000";
      when 17748 => pixel <= "000000";
      when 17749 => pixel <= "000000";
      when 17750 => pixel <= "000000";
      when 17751 => pixel <= "000000";
      when 17752 => pixel <= "000000";
      when 17753 => pixel <= "000000";
      when 17754 => pixel <= "000000";
      when 17755 => pixel <= "000000";
      when 17756 => pixel <= "000000";
      when 17757 => pixel <= "000000";
      when 17758 => pixel <= "000000";
      when 17759 => pixel <= "000000";
      when 17760 => pixel <= "000000";
      when 17761 => pixel <= "000000";
      when 17762 => pixel <= "000000";
      when 17763 => pixel <= "000000";
      when 17764 => pixel <= "000000";
      when 17765 => pixel <= "000000";
      when 17766 => pixel <= "000000";
      when 17767 => pixel <= "000000";
      when 17768 => pixel <= "000000";
      when 17769 => pixel <= "000000";
      when 17770 => pixel <= "000000";
      when 17771 => pixel <= "000000";
      when 17772 => pixel <= "000000";
      when 17773 => pixel <= "000000";
      when 17774 => pixel <= "000000";
      when 17775 => pixel <= "000000";
      when 17776 => pixel <= "000000";
      when 17777 => pixel <= "000000";
      when 17778 => pixel <= "000000";
      when 17779 => pixel <= "000000";
      when 17780 => pixel <= "000000";
      when 17781 => pixel <= "000000";
      when 17782 => pixel <= "000000";
      when 17783 => pixel <= "000000";
      when 17784 => pixel <= "000000";
      when 17785 => pixel <= "000000";
      when 17786 => pixel <= "000000";
      when 17787 => pixel <= "000000";
      when 17788 => pixel <= "000000";
      when 17789 => pixel <= "000000";
      when 17790 => pixel <= "000000";
      when 17791 => pixel <= "000000";
      when 17792 => pixel <= "000000";
      when 17793 => pixel <= "000000";
      when 17794 => pixel <= "000000";
      when 17795 => pixel <= "000000";
      when 17796 => pixel <= "000000";
      when 17797 => pixel <= "000000";
      when 17798 => pixel <= "000000";
      when 17799 => pixel <= "000000";
      when 17800 => pixel <= "000000";
      when 17801 => pixel <= "000000";
      when 17802 => pixel <= "000000";
      when 17803 => pixel <= "000000";
      when 17804 => pixel <= "000000";
      when 17805 => pixel <= "000000";
      when 17806 => pixel <= "000000";
      when 17807 => pixel <= "000000";
      when 17808 => pixel <= "000000";
      when 17809 => pixel <= "000000";
      when 17810 => pixel <= "000000";
      when 17811 => pixel <= "000000";
      when 17812 => pixel <= "000000";
      when 17813 => pixel <= "000000";
      when 17814 => pixel <= "000000";
      when 17815 => pixel <= "000000";
      when 17816 => pixel <= "000000";
      when 17817 => pixel <= "000000";
      when 17818 => pixel <= "000000";
      when 17819 => pixel <= "000000";
      when 17820 => pixel <= "000000";
      when 17821 => pixel <= "000000";
      when 17822 => pixel <= "000000";
      when 17823 => pixel <= "000000";
      when 17824 => pixel <= "000000";
      when 17825 => pixel <= "000000";
      when 17826 => pixel <= "000000";
      when 17827 => pixel <= "000000";
      when 17828 => pixel <= "000000";
      when 17829 => pixel <= "000000";
      when 17830 => pixel <= "000000";
      when 17831 => pixel <= "000000";
      when 17832 => pixel <= "000000";
      when 17833 => pixel <= "000000";
      when 17834 => pixel <= "000000";
      when 17835 => pixel <= "000000";
      when 17836 => pixel <= "000000";
      when 17837 => pixel <= "000000";
      when 17838 => pixel <= "000000";
      when 17839 => pixel <= "000000";
      when 17840 => pixel <= "000000";
      when 17841 => pixel <= "000000";
      when 17842 => pixel <= "000000";
      when 17843 => pixel <= "000000";
      when 17844 => pixel <= "000000";
      when 17845 => pixel <= "000000";
      when 17846 => pixel <= "000000";
      when 17847 => pixel <= "000000";
      when 17848 => pixel <= "000000";
      when 17849 => pixel <= "000000";
      when 17850 => pixel <= "000000";
      when 17851 => pixel <= "000000";
      when 17852 => pixel <= "000000";
      when 17853 => pixel <= "000000";
      when 17854 => pixel <= "000000";
      when 17855 => pixel <= "000000";
      when 17856 => pixel <= "000000";
      when 17857 => pixel <= "000000";
      when 17858 => pixel <= "000000";
      when 17859 => pixel <= "000000";
      when 17860 => pixel <= "000000";
      when 17861 => pixel <= "000000";
      when 17862 => pixel <= "000000";
      when 17863 => pixel <= "000000";
      when 17864 => pixel <= "000000";
      when 17865 => pixel <= "000000";
      when 17866 => pixel <= "000000";
      when 17867 => pixel <= "000000";
      when 17868 => pixel <= "000000";
      when 17869 => pixel <= "000000";
      when 17870 => pixel <= "000000";
      when 17871 => pixel <= "000000";
      when 17872 => pixel <= "000000";
      when 17873 => pixel <= "000000";
      when 17874 => pixel <= "000000";
      when 17875 => pixel <= "000000";
      when 17876 => pixel <= "000000";
      when 17877 => pixel <= "000000";
      when 17878 => pixel <= "000000";
      when 17879 => pixel <= "000000";
      when 17880 => pixel <= "000000";
      when 17881 => pixel <= "000000";
      when 17882 => pixel <= "000000";
      when 17883 => pixel <= "000000";
      when 17884 => pixel <= "000000";
      when 17885 => pixel <= "000000";
      when 17886 => pixel <= "000000";
      when 17887 => pixel <= "000000";
      when 17888 => pixel <= "000000";
      when 17889 => pixel <= "000000";
      when 17890 => pixel <= "000000";
      when 17891 => pixel <= "000000";
      when 17892 => pixel <= "000000";
      when 17893 => pixel <= "000000";
      when 17894 => pixel <= "000000";
      when 17895 => pixel <= "000000";
      when 17896 => pixel <= "000000";
      when 17897 => pixel <= "000000";
      when 17898 => pixel <= "000000";
      when 17899 => pixel <= "000000";
      when 17900 => pixel <= "000000";
      when 17901 => pixel <= "000000";
      when 17902 => pixel <= "000000";
      when 17903 => pixel <= "000000";
      when 17904 => pixel <= "000000";
      when 17905 => pixel <= "000000";
      when 17906 => pixel <= "000000";
      when 17907 => pixel <= "000000";
      when 17908 => pixel <= "000000";
      when 17909 => pixel <= "000000";
      when 17910 => pixel <= "000000";
      when 17911 => pixel <= "000000";
      when 17912 => pixel <= "000000";
      when 17913 => pixel <= "000000";
      when 17914 => pixel <= "000000";
      when 17915 => pixel <= "000000";
      when 17916 => pixel <= "000000";
      when 17917 => pixel <= "000000";
      when 17918 => pixel <= "000000";
      when 17919 => pixel <= "000000";
      when 17920 => pixel <= "000000";
      when 17921 => pixel <= "000000";
      when 17922 => pixel <= "000000";
      when 17923 => pixel <= "000000";
      when 17924 => pixel <= "000000";
      when 17925 => pixel <= "000000";
      when 17926 => pixel <= "000000";
      when 17927 => pixel <= "000000";
      when 17928 => pixel <= "000000";
      when 17929 => pixel <= "000000";
      when 17930 => pixel <= "000000";
      when 17931 => pixel <= "000000";
      when 17932 => pixel <= "000000";
      when 17933 => pixel <= "000000";
      when 17934 => pixel <= "000000";
      when 17935 => pixel <= "000000";
      when 17936 => pixel <= "000000";
      when 17937 => pixel <= "000000";
      when 17938 => pixel <= "000000";
      when 17939 => pixel <= "000000";
      when 17940 => pixel <= "000000";
      when 17941 => pixel <= "000000";
      when 17942 => pixel <= "000000";
      when 17943 => pixel <= "000000";
      when 17944 => pixel <= "000000";
      when 17945 => pixel <= "000000";
      when 17946 => pixel <= "000000";
      when 17947 => pixel <= "000000";
      when 17948 => pixel <= "000000";
      when 17949 => pixel <= "000000";
      when 17950 => pixel <= "000000";
      when 17951 => pixel <= "000000";
      when 17952 => pixel <= "000000";
      when 17953 => pixel <= "000000";
      when 17954 => pixel <= "000000";
      when 17955 => pixel <= "000000";
      when 17956 => pixel <= "000000";
      when 17957 => pixel <= "000000";
      when 17958 => pixel <= "000000";
      when 17959 => pixel <= "000000";
      when 17960 => pixel <= "000000";
      when 17961 => pixel <= "000000";
      when 17962 => pixel <= "000000";
      when 17963 => pixel <= "000000";
      when 17964 => pixel <= "000000";
      when 17965 => pixel <= "000000";
      when 17966 => pixel <= "000000";
      when 17967 => pixel <= "000000";
      when 17968 => pixel <= "000000";
      when 17969 => pixel <= "000000";
      when 17970 => pixel <= "000000";
      when 17971 => pixel <= "000000";
      when 17972 => pixel <= "000000";
      when 17973 => pixel <= "000000";
      when 17974 => pixel <= "000000";
      when 17975 => pixel <= "000000";
      when 17976 => pixel <= "000000";
      when 17977 => pixel <= "000000";
      when 17978 => pixel <= "000000";
      when 17979 => pixel <= "000000";
      when 17980 => pixel <= "000000";
      when 17981 => pixel <= "000000";
      when 17982 => pixel <= "000000";
      when 17983 => pixel <= "000000";
      when 17984 => pixel <= "000000";
      when 17985 => pixel <= "000000";
      when 17986 => pixel <= "000000";
      when 17987 => pixel <= "000000";
      when 17988 => pixel <= "000000";
      when 17989 => pixel <= "000000";
      when 17990 => pixel <= "000000";
      when 17991 => pixel <= "000000";
      when 17992 => pixel <= "000000";
      when 17993 => pixel <= "000000";
      when 17994 => pixel <= "000000";
      when 17995 => pixel <= "000000";
      when 17996 => pixel <= "000000";
      when 17997 => pixel <= "000000";
      when 17998 => pixel <= "000000";
      when 17999 => pixel <= "000000";
      when 18000 => pixel <= "000000";
      when 18001 => pixel <= "000000";
      when 18002 => pixel <= "000000";
      when 18003 => pixel <= "000000";
      when 18004 => pixel <= "000000";
      when 18005 => pixel <= "000000";
      when 18006 => pixel <= "000000";
      when 18007 => pixel <= "000000";
      when 18008 => pixel <= "000000";
      when 18009 => pixel <= "000000";
      when 18010 => pixel <= "000000";
      when 18011 => pixel <= "000000";
      when 18012 => pixel <= "000000";
      when 18013 => pixel <= "000000";
      when 18014 => pixel <= "000000";
      when 18015 => pixel <= "000000";
      when 18016 => pixel <= "000000";
      when 18017 => pixel <= "000000";
      when 18018 => pixel <= "000000";
      when 18019 => pixel <= "000000";
      when 18020 => pixel <= "000000";
      when 18021 => pixel <= "000000";
      when 18022 => pixel <= "000000";
      when 18023 => pixel <= "000000";
      when 18024 => pixel <= "000000";
      when 18025 => pixel <= "000000";
      when 18026 => pixel <= "000000";
      when 18027 => pixel <= "000000";
      when 18028 => pixel <= "000000";
      when 18029 => pixel <= "000000";
      when 18030 => pixel <= "000000";
      when 18031 => pixel <= "000000";
      when 18032 => pixel <= "000000";
      when 18033 => pixel <= "000000";
      when 18034 => pixel <= "000000";
      when 18035 => pixel <= "000000";
      when 18036 => pixel <= "000000";
      when 18037 => pixel <= "000000";
      when 18038 => pixel <= "000000";
      when 18039 => pixel <= "000000";
      when 18040 => pixel <= "000000";
      when 18041 => pixel <= "000000";
      when 18042 => pixel <= "000000";
      when 18043 => pixel <= "000000";
      when 18044 => pixel <= "000000";
      when 18045 => pixel <= "000000";
      when 18046 => pixel <= "000000";
      when 18047 => pixel <= "000000";
      when 18048 => pixel <= "000000";
      when 18049 => pixel <= "000000";
      when 18050 => pixel <= "000000";
      when 18051 => pixel <= "000000";
      when 18052 => pixel <= "000000";
      when 18053 => pixel <= "000000";
      when 18054 => pixel <= "000000";
      when 18055 => pixel <= "000000";
      when 18056 => pixel <= "000000";
      when 18057 => pixel <= "000000";
      when 18058 => pixel <= "000000";
      when 18059 => pixel <= "000000";
      when 18060 => pixel <= "000000";
      when 18061 => pixel <= "000000";
      when 18062 => pixel <= "000000";
      when 18063 => pixel <= "000000";
      when 18064 => pixel <= "000000";
      when 18065 => pixel <= "000000";
      when 18066 => pixel <= "000000";
      when 18067 => pixel <= "000000";
      when 18068 => pixel <= "000000";
      when 18069 => pixel <= "000000";
      when 18070 => pixel <= "000000";
      when 18071 => pixel <= "000000";
      when 18072 => pixel <= "000000";
      when 18073 => pixel <= "000000";
      when 18074 => pixel <= "000000";
      when 18075 => pixel <= "000000";
      when 18076 => pixel <= "000000";
      when 18077 => pixel <= "000000";
      when 18078 => pixel <= "000000";
      when 18079 => pixel <= "000000";
      when 18080 => pixel <= "000000";
      when 18081 => pixel <= "000000";
      when 18082 => pixel <= "000000";
      when 18083 => pixel <= "000000";
      when 18084 => pixel <= "000000";
      when 18085 => pixel <= "000000";
      when 18086 => pixel <= "000000";
      when 18087 => pixel <= "000000";
      when 18088 => pixel <= "000000";
      when 18089 => pixel <= "000000";
      when 18090 => pixel <= "000000";
      when 18091 => pixel <= "000000";
      when 18092 => pixel <= "000000";
      when 18093 => pixel <= "000000";
      when 18094 => pixel <= "000000";
      when 18095 => pixel <= "000000";
      when 18096 => pixel <= "000000";
      when 18097 => pixel <= "000000";
      when 18098 => pixel <= "000000";
      when 18099 => pixel <= "000000";
      when 18100 => pixel <= "000000";
      when 18101 => pixel <= "000000";
      when 18102 => pixel <= "000000";
      when 18103 => pixel <= "000000";
      when 18104 => pixel <= "000000";
      when 18105 => pixel <= "000000";
      when 18106 => pixel <= "000000";
      when 18107 => pixel <= "000000";
      when 18108 => pixel <= "000000";
      when 18109 => pixel <= "000000";
      when 18110 => pixel <= "000000";
      when 18111 => pixel <= "000000";
      when 18112 => pixel <= "000000";
      when 18113 => pixel <= "000000";
      when 18114 => pixel <= "000000";
      when 18115 => pixel <= "000000";
      when 18116 => pixel <= "000000";
      when 18117 => pixel <= "000000";
      when 18118 => pixel <= "000000";
      when 18119 => pixel <= "000000";
      when 18120 => pixel <= "000000";
      when 18121 => pixel <= "000000";
      when 18122 => pixel <= "000000";
      when 18123 => pixel <= "000000";
      when 18124 => pixel <= "000000";
      when 18125 => pixel <= "000000";
      when 18126 => pixel <= "000000";
      when 18127 => pixel <= "000000";
      when 18128 => pixel <= "000000";
      when 18129 => pixel <= "000000";
      when 18130 => pixel <= "000000";
      when 18131 => pixel <= "000000";
      when 18132 => pixel <= "000000";
      when 18133 => pixel <= "000000";
      when 18134 => pixel <= "000000";
      when 18135 => pixel <= "000000";
      when 18136 => pixel <= "000000";
      when 18137 => pixel <= "000000";
      when 18138 => pixel <= "000000";
      when 18139 => pixel <= "000000";
      when 18140 => pixel <= "000000";
      when 18141 => pixel <= "000000";
      when 18142 => pixel <= "000000";
      when 18143 => pixel <= "000000";
      when 18144 => pixel <= "000000";
      when 18145 => pixel <= "000000";
      when 18146 => pixel <= "000000";
      when 18147 => pixel <= "000000";
      when 18148 => pixel <= "000000";
      when 18149 => pixel <= "000000";
      when 18150 => pixel <= "000000";
      when 18151 => pixel <= "000000";
      when 18152 => pixel <= "000000";
      when 18153 => pixel <= "000000";
      when 18154 => pixel <= "000000";
      when 18155 => pixel <= "000000";
      when 18156 => pixel <= "000000";
      when 18157 => pixel <= "000000";
      when 18158 => pixel <= "000000";
      when 18159 => pixel <= "000000";
      when 18160 => pixel <= "000000";
      when 18161 => pixel <= "000000";
      when 18162 => pixel <= "000000";
      when 18163 => pixel <= "000000";
      when 18164 => pixel <= "000000";
      when 18165 => pixel <= "000000";
      when 18166 => pixel <= "000000";
      when 18167 => pixel <= "000000";
      when 18168 => pixel <= "000000";
      when 18169 => pixel <= "000000";
      when 18170 => pixel <= "000000";
      when 18171 => pixel <= "000000";
      when 18172 => pixel <= "000000";
      when 18173 => pixel <= "000000";
      when 18174 => pixel <= "000000";
      when 18175 => pixel <= "000000";
      when 18176 => pixel <= "000000";
      when 18177 => pixel <= "000000";
      when 18178 => pixel <= "000000";
      when 18179 => pixel <= "000000";
      when 18180 => pixel <= "000000";
      when 18181 => pixel <= "000000";
      when 18182 => pixel <= "000000";
      when 18183 => pixel <= "000000";
      when 18184 => pixel <= "000000";
      when 18185 => pixel <= "000000";
      when 18186 => pixel <= "000000";
      when 18187 => pixel <= "000000";
      when 18188 => pixel <= "000000";
      when 18189 => pixel <= "000000";
      when 18190 => pixel <= "000000";
      when 18191 => pixel <= "000000";
      when 18192 => pixel <= "000000";
      when 18193 => pixel <= "000000";
      when 18194 => pixel <= "000000";
      when 18195 => pixel <= "000000";
      when 18196 => pixel <= "000000";
      when 18197 => pixel <= "000000";
      when 18198 => pixel <= "000000";
      when 18199 => pixel <= "000000";
      when 18200 => pixel <= "000000";
      when 18201 => pixel <= "000000";
      when 18202 => pixel <= "000000";
      when 18203 => pixel <= "000000";
      when 18204 => pixel <= "000000";
      when 18205 => pixel <= "000000";
      when 18206 => pixel <= "000000";
      when 18207 => pixel <= "000000";
      when 18208 => pixel <= "000000";
      when 18209 => pixel <= "000000";
      when 18210 => pixel <= "000000";
      when 18211 => pixel <= "000000";
      when 18212 => pixel <= "000000";
      when 18213 => pixel <= "000000";
      when 18214 => pixel <= "000000";
      when 18215 => pixel <= "000000";
      when 18216 => pixel <= "000000";
      when 18217 => pixel <= "000000";
      when 18218 => pixel <= "000000";
      when 18219 => pixel <= "000000";
      when 18220 => pixel <= "000000";
      when 18221 => pixel <= "000000";
      when 18222 => pixel <= "000000";
      when 18223 => pixel <= "000000";
      when 18224 => pixel <= "000000";
      when 18225 => pixel <= "000000";
      when 18226 => pixel <= "000000";
      when 18227 => pixel <= "000000";
      when 18228 => pixel <= "000000";
      when 18229 => pixel <= "000000";
      when 18230 => pixel <= "000000";
      when 18231 => pixel <= "000000";
      when 18232 => pixel <= "000000";
      when 18233 => pixel <= "000000";
      when 18234 => pixel <= "000000";
      when 18235 => pixel <= "000000";
      when 18236 => pixel <= "000000";
      when 18237 => pixel <= "000000";
      when 18238 => pixel <= "000000";
      when 18239 => pixel <= "000000";
      when 18240 => pixel <= "000000";
      when 18241 => pixel <= "000000";
      when 18242 => pixel <= "000000";
      when 18243 => pixel <= "000000";
      when 18244 => pixel <= "000000";
      when 18245 => pixel <= "000000";
      when 18246 => pixel <= "000000";
      when 18247 => pixel <= "000000";
      when 18248 => pixel <= "000000";
      when 18249 => pixel <= "000000";
      when 18250 => pixel <= "000000";
      when 18251 => pixel <= "000000";
      when 18252 => pixel <= "000000";
      when 18253 => pixel <= "000000";
      when 18254 => pixel <= "000000";
      when 18255 => pixel <= "000000";
      when 18256 => pixel <= "000000";
      when 18257 => pixel <= "000000";
      when 18258 => pixel <= "000000";
      when 18259 => pixel <= "000000";
      when 18260 => pixel <= "000000";
      when 18261 => pixel <= "000000";
      when 18262 => pixel <= "000000";
      when 18263 => pixel <= "000000";
      when 18264 => pixel <= "000000";
      when 18265 => pixel <= "000000";
      when 18266 => pixel <= "000000";
      when 18267 => pixel <= "000000";
      when 18268 => pixel <= "000000";
      when 18269 => pixel <= "000000";
      when 18270 => pixel <= "000000";
      when 18271 => pixel <= "000000";
      when 18272 => pixel <= "000000";
      when 18273 => pixel <= "000000";
      when 18274 => pixel <= "000000";
      when 18275 => pixel <= "000000";
      when 18276 => pixel <= "000000";
      when 18277 => pixel <= "000000";
      when 18278 => pixel <= "000000";
      when 18279 => pixel <= "000000";
      when 18280 => pixel <= "000000";
      when 18281 => pixel <= "000000";
      when 18282 => pixel <= "000000";
      when 18283 => pixel <= "000000";
      when 18284 => pixel <= "000000";
      when 18285 => pixel <= "000000";
      when 18286 => pixel <= "000000";
      when 18287 => pixel <= "000000";
      when 18288 => pixel <= "000000";
      when 18289 => pixel <= "000000";
      when 18290 => pixel <= "000000";
      when 18291 => pixel <= "000000";
      when 18292 => pixel <= "000000";
      when 18293 => pixel <= "000000";
      when 18294 => pixel <= "000000";
      when 18295 => pixel <= "000000";
      when 18296 => pixel <= "000000";
      when 18297 => pixel <= "000000";
      when 18298 => pixel <= "000000";
      when 18299 => pixel <= "000000";
      when 18300 => pixel <= "000000";
      when 18301 => pixel <= "000000";
      when 18302 => pixel <= "000000";
      when 18303 => pixel <= "000000";
      when 18304 => pixel <= "000000";
      when 18305 => pixel <= "000000";
      when 18306 => pixel <= "000000";
      when 18307 => pixel <= "000000";
      when 18308 => pixel <= "000000";
      when 18309 => pixel <= "000000";
      when 18310 => pixel <= "000000";
      when 18311 => pixel <= "000000";
      when 18312 => pixel <= "000000";
      when 18313 => pixel <= "000000";
      when 18314 => pixel <= "000000";
      when 18315 => pixel <= "000000";
      when 18316 => pixel <= "000000";
      when 18317 => pixel <= "000000";
      when 18318 => pixel <= "000000";
      when 18319 => pixel <= "000000";
      when 18320 => pixel <= "000000";
      when 18321 => pixel <= "000000";
      when 18322 => pixel <= "000000";
      when 18323 => pixel <= "000000";
      when 18324 => pixel <= "000000";
      when 18325 => pixel <= "000000";
      when 18326 => pixel <= "000000";
      when 18327 => pixel <= "000000";
      when 18328 => pixel <= "000000";
      when 18329 => pixel <= "000000";
      when 18330 => pixel <= "000000";
      when 18331 => pixel <= "000000";
      when 18332 => pixel <= "000000";
      when 18333 => pixel <= "000000";
      when 18334 => pixel <= "000000";
      when 18335 => pixel <= "000000";
      when 18336 => pixel <= "000000";
      when 18337 => pixel <= "000000";
      when 18338 => pixel <= "000000";
      when 18339 => pixel <= "000000";
      when 18340 => pixel <= "000000";
      when 18341 => pixel <= "000000";
      when 18342 => pixel <= "000000";
      when 18343 => pixel <= "000000";
      when 18344 => pixel <= "000000";
      when 18345 => pixel <= "000000";
      when 18346 => pixel <= "000000";
      when 18347 => pixel <= "000000";
      when 18348 => pixel <= "000000";
      when 18349 => pixel <= "000000";
      when 18350 => pixel <= "000000";
      when 18351 => pixel <= "000000";
      when 18352 => pixel <= "000000";
      when 18353 => pixel <= "000000";
      when 18354 => pixel <= "000000";
      when 18355 => pixel <= "000000";
      when 18356 => pixel <= "000000";
      when 18357 => pixel <= "000000";
      when 18358 => pixel <= "000000";
      when 18359 => pixel <= "000000";
      when 18360 => pixel <= "000000";
      when 18361 => pixel <= "000000";
      when 18362 => pixel <= "000000";
      when 18363 => pixel <= "000000";
      when 18364 => pixel <= "000000";
      when 18365 => pixel <= "000000";
      when 18366 => pixel <= "000000";
      when 18367 => pixel <= "000000";
      when 18368 => pixel <= "000000";
      when 18369 => pixel <= "000000";
      when 18370 => pixel <= "000000";
      when 18371 => pixel <= "000000";
      when 18372 => pixel <= "000000";
      when 18373 => pixel <= "000000";
      when 18374 => pixel <= "000000";
      when 18375 => pixel <= "000000";
      when 18376 => pixel <= "000000";
      when 18377 => pixel <= "000000";
      when 18378 => pixel <= "000000";
      when 18379 => pixel <= "000000";
      when 18380 => pixel <= "000000";
      when 18381 => pixel <= "000000";
      when 18382 => pixel <= "000000";
      when 18383 => pixel <= "000000";
      when 18384 => pixel <= "000000";
      when 18385 => pixel <= "000000";
      when 18386 => pixel <= "000000";
      when 18387 => pixel <= "000000";
      when 18388 => pixel <= "000000";
      when 18389 => pixel <= "000000";
      when 18390 => pixel <= "000000";
      when 18391 => pixel <= "000000";
      when 18392 => pixel <= "000000";
      when 18393 => pixel <= "000000";
      when 18394 => pixel <= "000000";
      when 18395 => pixel <= "000000";
      when 18396 => pixel <= "000000";
      when 18397 => pixel <= "000000";
      when 18398 => pixel <= "000000";
      when 18399 => pixel <= "000000";
      when 18400 => pixel <= "000000";
      when 18401 => pixel <= "000000";
      when 18402 => pixel <= "000000";
      when 18403 => pixel <= "000000";
      when 18404 => pixel <= "000000";
      when 18405 => pixel <= "000000";
      when 18406 => pixel <= "000000";
      when 18407 => pixel <= "000000";
      when 18408 => pixel <= "000000";
      when 18409 => pixel <= "000000";
      when 18410 => pixel <= "000000";
      when 18411 => pixel <= "000000";
      when 18412 => pixel <= "000000";
      when 18413 => pixel <= "000000";
      when 18414 => pixel <= "000000";
      when 18415 => pixel <= "000000";
      when 18416 => pixel <= "000000";
      when 18417 => pixel <= "000000";
      when 18418 => pixel <= "000000";
      when 18419 => pixel <= "000000";
      when 18420 => pixel <= "000000";
      when 18421 => pixel <= "000000";
      when 18422 => pixel <= "000000";
      when 18423 => pixel <= "000000";
      when 18424 => pixel <= "000000";
      when 18425 => pixel <= "000000";
      when 18426 => pixel <= "000000";
      when 18427 => pixel <= "000000";
      when 18428 => pixel <= "000000";
      when 18429 => pixel <= "000000";
      when 18430 => pixel <= "000000";
      when 18431 => pixel <= "000000";
      when 18432 => pixel <= "000000";
      when 18433 => pixel <= "000000";
      when 18434 => pixel <= "000000";
      when 18435 => pixel <= "000000";
      when 18436 => pixel <= "000000";
      when 18437 => pixel <= "000000";
      when 18438 => pixel <= "000000";
      when 18439 => pixel <= "000000";
      when 18440 => pixel <= "000000";
      when 18441 => pixel <= "000000";
      when 18442 => pixel <= "000000";
      when 18443 => pixel <= "000000";
      when 18444 => pixel <= "000000";
      when 18445 => pixel <= "000000";
      when 18446 => pixel <= "000000";
      when 18447 => pixel <= "000000";
      when 18448 => pixel <= "000000";
      when 18449 => pixel <= "000000";
      when 18450 => pixel <= "000000";
      when 18451 => pixel <= "000000";
      when 18452 => pixel <= "000000";
      when 18453 => pixel <= "000000";
      when 18454 => pixel <= "000000";
      when 18455 => pixel <= "000000";
      when 18456 => pixel <= "000000";
      when 18457 => pixel <= "000000";
      when 18458 => pixel <= "000000";
      when 18459 => pixel <= "000000";
      when 18460 => pixel <= "000000";
      when 18461 => pixel <= "000000";
      when 18462 => pixel <= "000000";
      when 18463 => pixel <= "000000";
      when 18464 => pixel <= "000000";
      when 18465 => pixel <= "000000";
      when 18466 => pixel <= "000000";
      when 18467 => pixel <= "000000";
      when 18468 => pixel <= "000000";
      when 18469 => pixel <= "000000";
      when 18470 => pixel <= "000000";
      when 18471 => pixel <= "000000";
      when 18472 => pixel <= "000000";
      when 18473 => pixel <= "000000";
      when 18474 => pixel <= "000000";
      when 18475 => pixel <= "000000";
      when 18476 => pixel <= "000000";
      when 18477 => pixel <= "000000";
      when 18478 => pixel <= "000000";
      when 18479 => pixel <= "000000";
      when 18480 => pixel <= "000000";
      when 18481 => pixel <= "000000";
      when 18482 => pixel <= "000000";
      when 18483 => pixel <= "000000";
      when 18484 => pixel <= "000000";
      when 18485 => pixel <= "000000";
      when 18486 => pixel <= "000000";
      when 18487 => pixel <= "000000";
      when 18488 => pixel <= "000000";
      when 18489 => pixel <= "000000";
      when 18490 => pixel <= "000000";
      when 18491 => pixel <= "000000";
      when 18492 => pixel <= "000000";
      when 18493 => pixel <= "000000";
      when 18494 => pixel <= "000000";
      when 18495 => pixel <= "000000";
      when 18496 => pixel <= "000000";
      when 18497 => pixel <= "000000";
      when 18498 => pixel <= "000000";
      when 18499 => pixel <= "000000";
      when 18500 => pixel <= "000000";
      when 18501 => pixel <= "000000";
      when 18502 => pixel <= "000000";
      when 18503 => pixel <= "000000";
      when 18504 => pixel <= "000000";
      when 18505 => pixel <= "000000";
      when 18506 => pixel <= "000000";
      when 18507 => pixel <= "000000";
      when 18508 => pixel <= "000000";
      when 18509 => pixel <= "000000";
      when 18510 => pixel <= "000000";
      when 18511 => pixel <= "000000";
      when 18512 => pixel <= "000000";
      when 18513 => pixel <= "000000";
      when 18514 => pixel <= "000000";
      when 18515 => pixel <= "000000";
      when 18516 => pixel <= "000000";
      when 18517 => pixel <= "000000";
      when 18518 => pixel <= "000000";
      when 18519 => pixel <= "000000";
      when 18520 => pixel <= "000000";
      when 18521 => pixel <= "000000";
      when 18522 => pixel <= "000000";
      when 18523 => pixel <= "000000";
      when 18524 => pixel <= "000000";
      when 18525 => pixel <= "000000";
      when 18526 => pixel <= "000000";
      when 18527 => pixel <= "000000";
      when 18528 => pixel <= "000000";
      when 18529 => pixel <= "000000";
      when 18530 => pixel <= "000000";
      when 18531 => pixel <= "000000";
      when 18532 => pixel <= "000000";
      when 18533 => pixel <= "000000";
      when 18534 => pixel <= "000000";
      when 18535 => pixel <= "000000";
      when 18536 => pixel <= "000000";
      when 18537 => pixel <= "000000";
      when 18538 => pixel <= "000000";
      when 18539 => pixel <= "000000";
      when 18540 => pixel <= "000000";
      when 18541 => pixel <= "000000";
      when 18542 => pixel <= "000000";
      when 18543 => pixel <= "000000";
      when 18544 => pixel <= "000000";
      when 18545 => pixel <= "000000";
      when 18546 => pixel <= "000000";
      when 18547 => pixel <= "000000";
      when 18548 => pixel <= "000000";
      when 18549 => pixel <= "000000";
      when 18550 => pixel <= "000000";
      when 18551 => pixel <= "000000";
      when 18552 => pixel <= "000000";
      when 18553 => pixel <= "000000";
      when 18554 => pixel <= "000000";
      when 18555 => pixel <= "000000";
      when 18556 => pixel <= "000000";
      when 18557 => pixel <= "000000";
      when 18558 => pixel <= "000000";
      when 18559 => pixel <= "000000";
      when 18560 => pixel <= "000000";
      when 18561 => pixel <= "000000";
      when 18562 => pixel <= "000000";
      when 18563 => pixel <= "000000";
      when 18564 => pixel <= "000000";
      when 18565 => pixel <= "000000";
      when 18566 => pixel <= "000000";
      when 18567 => pixel <= "000000";
      when 18568 => pixel <= "000000";
      when 18569 => pixel <= "000000";
      when 18570 => pixel <= "000000";
      when 18571 => pixel <= "000000";
      when 18572 => pixel <= "000000";
      when 18573 => pixel <= "000000";
      when 18574 => pixel <= "000000";
      when 18575 => pixel <= "000000";
      when 18576 => pixel <= "000000";
      when 18577 => pixel <= "000000";
      when 18578 => pixel <= "000000";
      when 18579 => pixel <= "000000";
      when 18580 => pixel <= "000000";
      when 18581 => pixel <= "000000";
      when 18582 => pixel <= "000000";
      when 18583 => pixel <= "000000";
      when 18584 => pixel <= "000000";
      when 18585 => pixel <= "000000";
      when 18586 => pixel <= "000000";
      when 18587 => pixel <= "000000";
      when 18588 => pixel <= "000000";
      when 18589 => pixel <= "000000";
      when 18590 => pixel <= "000000";
      when 18591 => pixel <= "000000";
      when 18592 => pixel <= "000000";
      when 18593 => pixel <= "000000";
      when 18594 => pixel <= "000000";
      when 18595 => pixel <= "000000";
      when 18596 => pixel <= "000000";
      when 18597 => pixel <= "000000";
      when 18598 => pixel <= "000000";
      when 18599 => pixel <= "000000";
      when 18600 => pixel <= "000000";
      when 18601 => pixel <= "000000";
      when 18602 => pixel <= "000000";
      when 18603 => pixel <= "000000";
      when 18604 => pixel <= "000000";
      when 18605 => pixel <= "000000";
      when 18606 => pixel <= "000000";
      when 18607 => pixel <= "000000";
      when 18608 => pixel <= "000000";
      when 18609 => pixel <= "000000";
      when 18610 => pixel <= "000000";
      when 18611 => pixel <= "000000";
      when 18612 => pixel <= "000000";
      when 18613 => pixel <= "000000";
      when 18614 => pixel <= "000000";
      when 18615 => pixel <= "000000";
      when 18616 => pixel <= "000000";
      when 18617 => pixel <= "000000";
      when 18618 => pixel <= "000000";
      when 18619 => pixel <= "000000";
      when 18620 => pixel <= "000000";
      when 18621 => pixel <= "000000";
      when 18622 => pixel <= "000000";
      when 18623 => pixel <= "000000";
      when 18624 => pixel <= "000000";
      when 18625 => pixel <= "000000";
      when 18626 => pixel <= "000000";
      when 18627 => pixel <= "000000";
      when 18628 => pixel <= "000000";
      when 18629 => pixel <= "000000";
      when 18630 => pixel <= "000000";
      when 18631 => pixel <= "000000";
      when 18632 => pixel <= "000000";
      when 18633 => pixel <= "000000";
      when 18634 => pixel <= "000000";
      when 18635 => pixel <= "000000";
      when 18636 => pixel <= "000000";
      when 18637 => pixel <= "000000";
      when 18638 => pixel <= "000000";
      when 18639 => pixel <= "000000";
      when 18640 => pixel <= "000000";
      when 18641 => pixel <= "000000";
      when 18642 => pixel <= "000000";
      when 18643 => pixel <= "000000";
      when 18644 => pixel <= "000000";
      when 18645 => pixel <= "000000";
      when 18646 => pixel <= "000000";
      when 18647 => pixel <= "000000";
      when 18648 => pixel <= "000000";
      when 18649 => pixel <= "000000";
      when 18650 => pixel <= "000000";
      when 18651 => pixel <= "000000";
      when 18652 => pixel <= "000000";
      when 18653 => pixel <= "000000";
      when 18654 => pixel <= "000000";
      when 18655 => pixel <= "000000";
      when 18656 => pixel <= "000000";
      when 18657 => pixel <= "000000";
      when 18658 => pixel <= "000000";
      when 18659 => pixel <= "000000";
      when 18660 => pixel <= "000000";
      when 18661 => pixel <= "000000";
      when 18662 => pixel <= "000000";
      when 18663 => pixel <= "000000";
      when 18664 => pixel <= "000000";
      when 18665 => pixel <= "000000";
      when 18666 => pixel <= "000000";
      when 18667 => pixel <= "000000";
      when 18668 => pixel <= "000000";
      when 18669 => pixel <= "000000";
      when 18670 => pixel <= "000000";
      when 18671 => pixel <= "000000";
      when 18672 => pixel <= "000000";
      when 18673 => pixel <= "000000";
      when 18674 => pixel <= "000000";
      when 18675 => pixel <= "000000";
      when 18676 => pixel <= "000000";
      when 18677 => pixel <= "000000";
      when 18678 => pixel <= "000000";
      when 18679 => pixel <= "000000";
      when 18680 => pixel <= "000000";
      when 18681 => pixel <= "000000";
      when 18682 => pixel <= "000000";
      when 18683 => pixel <= "000000";
      when 18684 => pixel <= "000000";
      when 18685 => pixel <= "000000";
      when 18686 => pixel <= "000000";
      when 18687 => pixel <= "000000";
      when 18688 => pixel <= "000000";
      when 18689 => pixel <= "000000";
      when 18690 => pixel <= "000000";
      when 18691 => pixel <= "000000";
      when 18692 => pixel <= "000000";
      when 18693 => pixel <= "000000";
      when 18694 => pixel <= "000000";
      when 18695 => pixel <= "000000";
      when 18696 => pixel <= "000000";
      when 18697 => pixel <= "000000";
      when 18698 => pixel <= "000000";
      when 18699 => pixel <= "000000";
      when 18700 => pixel <= "000000";
      when 18701 => pixel <= "000000";
      when 18702 => pixel <= "000000";
      when 18703 => pixel <= "000000";
      when 18704 => pixel <= "000000";
      when 18705 => pixel <= "000000";
      when 18706 => pixel <= "000000";
      when 18707 => pixel <= "000000";
      when 18708 => pixel <= "000000";
      when 18709 => pixel <= "000000";
      when 18710 => pixel <= "000000";
      when 18711 => pixel <= "000000";
      when 18712 => pixel <= "000000";
      when 18713 => pixel <= "000000";
      when 18714 => pixel <= "000000";
      when 18715 => pixel <= "000000";
      when 18716 => pixel <= "000000";
      when 18717 => pixel <= "000000";
      when 18718 => pixel <= "000000";
      when 18719 => pixel <= "000000";
      when 18720 => pixel <= "000000";
      when 18721 => pixel <= "000000";
      when 18722 => pixel <= "000000";
      when 18723 => pixel <= "000000";
      when 18724 => pixel <= "000000";
      when 18725 => pixel <= "000000";
      when 18726 => pixel <= "000000";
      when 18727 => pixel <= "000000";
      when 18728 => pixel <= "000000";
      when 18729 => pixel <= "000000";
      when 18730 => pixel <= "000000";
      when 18731 => pixel <= "000000";
      when 18732 => pixel <= "000000";
      when 18733 => pixel <= "000000";
      when 18734 => pixel <= "000000";
      when 18735 => pixel <= "000000";
      when 18736 => pixel <= "000000";
      when 18737 => pixel <= "000000";
      when 18738 => pixel <= "000000";
      when 18739 => pixel <= "000000";
      when 18740 => pixel <= "000000";
      when 18741 => pixel <= "000000";
      when 18742 => pixel <= "000000";
      when 18743 => pixel <= "000000";
      when 18744 => pixel <= "000000";
      when 18745 => pixel <= "000000";
      when 18746 => pixel <= "000000";
      when 18747 => pixel <= "000000";
      when 18748 => pixel <= "000000";
      when 18749 => pixel <= "000000";
      when 18750 => pixel <= "000000";
      when 18751 => pixel <= "000000";
      when 18752 => pixel <= "000000";
      when 18753 => pixel <= "000000";
      when 18754 => pixel <= "000000";
      when 18755 => pixel <= "000000";
      when 18756 => pixel <= "000000";
      when 18757 => pixel <= "000000";
      when 18758 => pixel <= "000000";
      when 18759 => pixel <= "000000";
      when 18760 => pixel <= "000000";
      when 18761 => pixel <= "000000";
      when 18762 => pixel <= "000000";
      when 18763 => pixel <= "000000";
      when 18764 => pixel <= "000000";
      when 18765 => pixel <= "000000";
      when 18766 => pixel <= "000000";
      when 18767 => pixel <= "000000";
      when 18768 => pixel <= "000000";
      when 18769 => pixel <= "000000";
      when 18770 => pixel <= "000000";
      when 18771 => pixel <= "000000";
      when 18772 => pixel <= "000000";
      when 18773 => pixel <= "000000";
      when 18774 => pixel <= "000000";
      when 18775 => pixel <= "000000";
      when 18776 => pixel <= "000000";
      when 18777 => pixel <= "000000";
      when 18778 => pixel <= "000000";
      when 18779 => pixel <= "000000";
      when 18780 => pixel <= "000000";
      when 18781 => pixel <= "000000";
      when 18782 => pixel <= "000000";
      when 18783 => pixel <= "000000";
      when 18784 => pixel <= "000000";
      when 18785 => pixel <= "000000";
      when 18786 => pixel <= "000000";
      when 18787 => pixel <= "000000";
      when 18788 => pixel <= "000000";
      when 18789 => pixel <= "000000";
      when 18790 => pixel <= "000000";
      when 18791 => pixel <= "000000";
      when 18792 => pixel <= "000000";
      when 18793 => pixel <= "000000";
      when 18794 => pixel <= "000000";
      when 18795 => pixel <= "000000";
      when 18796 => pixel <= "000000";
      when 18797 => pixel <= "000000";
      when 18798 => pixel <= "000000";
      when 18799 => pixel <= "000000";
      when 18800 => pixel <= "000000";
      when 18801 => pixel <= "000000";
      when 18802 => pixel <= "000000";
      when 18803 => pixel <= "000000";
      when 18804 => pixel <= "000000";
      when 18805 => pixel <= "000000";
      when 18806 => pixel <= "000000";
      when 18807 => pixel <= "000000";
      when 18808 => pixel <= "000000";
      when 18809 => pixel <= "000000";
      when 18810 => pixel <= "000000";
      when 18811 => pixel <= "000000";
      when 18812 => pixel <= "000000";
      when 18813 => pixel <= "000000";
      when 18814 => pixel <= "000000";
      when 18815 => pixel <= "000000";
      when 18816 => pixel <= "000000";
      when 18817 => pixel <= "000000";
      when 18818 => pixel <= "000000";
      when 18819 => pixel <= "000000";
      when 18820 => pixel <= "000000";
      when 18821 => pixel <= "000000";
      when 18822 => pixel <= "000000";
      when 18823 => pixel <= "000000";
      when 18824 => pixel <= "000000";
      when 18825 => pixel <= "000000";
      when 18826 => pixel <= "000000";
      when 18827 => pixel <= "000000";
      when 18828 => pixel <= "000000";
      when 18829 => pixel <= "000000";
      when 18830 => pixel <= "000000";
      when 18831 => pixel <= "000000";
      when 18832 => pixel <= "000000";
      when 18833 => pixel <= "000000";
      when 18834 => pixel <= "000000";
      when 18835 => pixel <= "000000";
      when 18836 => pixel <= "000000";
      when 18837 => pixel <= "000000";
      when 18838 => pixel <= "000000";
      when 18839 => pixel <= "000000";
      when 18840 => pixel <= "000000";
      when 18841 => pixel <= "000000";
      when 18842 => pixel <= "000000";
      when 18843 => pixel <= "000000";
      when 18844 => pixel <= "000000";
      when 18845 => pixel <= "000000";
      when 18846 => pixel <= "000000";
      when 18847 => pixel <= "000000";
      when 18848 => pixel <= "000000";
      when 18849 => pixel <= "000000";
      when 18850 => pixel <= "000000";
      when 18851 => pixel <= "000000";
      when 18852 => pixel <= "000000";
      when 18853 => pixel <= "000000";
      when 18854 => pixel <= "000000";
      when 18855 => pixel <= "000000";
      when 18856 => pixel <= "000000";
      when 18857 => pixel <= "000000";
      when 18858 => pixel <= "000000";
      when 18859 => pixel <= "000000";
      when 18860 => pixel <= "000000";
      when 18861 => pixel <= "000000";
      when 18862 => pixel <= "000000";
      when 18863 => pixel <= "000000";
      when 18864 => pixel <= "000000";
      when 18865 => pixel <= "000000";
      when 18866 => pixel <= "000000";
      when 18867 => pixel <= "000000";
      when 18868 => pixel <= "000000";
      when 18869 => pixel <= "000000";
      when 18870 => pixel <= "000000";
      when 18871 => pixel <= "000000";
      when 18872 => pixel <= "000000";
      when 18873 => pixel <= "000000";
      when 18874 => pixel <= "000000";
      when 18875 => pixel <= "000000";
      when 18876 => pixel <= "000000";
      when 18877 => pixel <= "000000";
      when 18878 => pixel <= "000000";
      when 18879 => pixel <= "000000";
      when 18880 => pixel <= "000000";
      when 18881 => pixel <= "000000";
      when 18882 => pixel <= "000000";
      when 18883 => pixel <= "000000";
      when 18884 => pixel <= "000000";
      when 18885 => pixel <= "000000";
      when 18886 => pixel <= "000000";
      when 18887 => pixel <= "000000";
      when 18888 => pixel <= "000000";
      when 18889 => pixel <= "000000";
      when 18890 => pixel <= "000000";
      when 18891 => pixel <= "000000";
      when 18892 => pixel <= "000000";
      when 18893 => pixel <= "000000";
      when 18894 => pixel <= "000000";
      when 18895 => pixel <= "000000";
      when 18896 => pixel <= "000000";
      when 18897 => pixel <= "000000";
      when 18898 => pixel <= "000000";
      when 18899 => pixel <= "000000";
      when 18900 => pixel <= "000000";
      when 18901 => pixel <= "000000";
      when 18902 => pixel <= "000000";
      when 18903 => pixel <= "000000";
      when 18904 => pixel <= "000000";
      when 18905 => pixel <= "000000";
      when 18906 => pixel <= "000000";
      when 18907 => pixel <= "000000";
      when 18908 => pixel <= "000000";
      when 18909 => pixel <= "000000";
      when 18910 => pixel <= "000000";
      when 18911 => pixel <= "000000";
      when 18912 => pixel <= "000000";
      when 18913 => pixel <= "000000";
      when 18914 => pixel <= "000000";
      when 18915 => pixel <= "000000";
      when 18916 => pixel <= "000000";
      when 18917 => pixel <= "000000";
      when 18918 => pixel <= "000000";
      when 18919 => pixel <= "000000";
      when 18920 => pixel <= "000000";
      when 18921 => pixel <= "000000";
      when 18922 => pixel <= "000000";
      when 18923 => pixel <= "000000";
      when 18924 => pixel <= "000000";
      when 18925 => pixel <= "000000";
      when 18926 => pixel <= "000000";
      when 18927 => pixel <= "000000";
      when 18928 => pixel <= "000000";
      when 18929 => pixel <= "000000";
      when 18930 => pixel <= "000000";
      when 18931 => pixel <= "000000";
      when 18932 => pixel <= "000000";
      when 18933 => pixel <= "000000";
      when 18934 => pixel <= "000000";
      when 18935 => pixel <= "000000";
      when 18936 => pixel <= "000000";
      when 18937 => pixel <= "000000";
      when 18938 => pixel <= "000000";
      when 18939 => pixel <= "000000";
      when 18940 => pixel <= "000000";
      when 18941 => pixel <= "000000";
      when 18942 => pixel <= "000000";
      when 18943 => pixel <= "000000";
      when 18944 => pixel <= "000000";
      when 18945 => pixel <= "000000";
      when 18946 => pixel <= "000000";
      when 18947 => pixel <= "000000";
      when 18948 => pixel <= "000000";
      when 18949 => pixel <= "000000";
      when 18950 => pixel <= "000000";
      when 18951 => pixel <= "000000";
      when 18952 => pixel <= "000000";
      when 18953 => pixel <= "000000";
      when 18954 => pixel <= "000000";
      when 18955 => pixel <= "000000";
      when 18956 => pixel <= "000000";
      when 18957 => pixel <= "000000";
      when 18958 => pixel <= "000000";
      when 18959 => pixel <= "000000";
      when 18960 => pixel <= "000000";
      when 18961 => pixel <= "000000";
      when 18962 => pixel <= "000000";
      when 18963 => pixel <= "000000";
      when 18964 => pixel <= "000000";
      when 18965 => pixel <= "000000";
      when 18966 => pixel <= "000000";
      when 18967 => pixel <= "000000";
      when 18968 => pixel <= "000000";
      when 18969 => pixel <= "000000";
      when 18970 => pixel <= "000000";
      when 18971 => pixel <= "000000";
      when 18972 => pixel <= "000000";
      when 18973 => pixel <= "000000";
      when 18974 => pixel <= "000000";
      when 18975 => pixel <= "000000";
      when 18976 => pixel <= "000000";
      when 18977 => pixel <= "000000";
      when 18978 => pixel <= "000000";
      when 18979 => pixel <= "000000";
      when 18980 => pixel <= "000000";
      when 18981 => pixel <= "000000";
      when 18982 => pixel <= "000000";
      when 18983 => pixel <= "000000";
      when 18984 => pixel <= "000000";
      when 18985 => pixel <= "000000";
      when 18986 => pixel <= "000000";
      when 18987 => pixel <= "000000";
      when 18988 => pixel <= "000000";
      when 18989 => pixel <= "000000";
      when 18990 => pixel <= "000000";
      when 18991 => pixel <= "000000";
      when 18992 => pixel <= "000000";
      when 18993 => pixel <= "000000";
      when 18994 => pixel <= "000000";
      when 18995 => pixel <= "000000";
      when 18996 => pixel <= "000000";
      when 18997 => pixel <= "000000";
      when 18998 => pixel <= "000000";
      when 18999 => pixel <= "000000";
      when 19000 => pixel <= "000000";
      when 19001 => pixel <= "000000";
      when 19002 => pixel <= "000000";
      when 19003 => pixel <= "000000";
      when 19004 => pixel <= "000000";
      when 19005 => pixel <= "000000";
      when 19006 => pixel <= "000000";
      when 19007 => pixel <= "000000";
      when 19008 => pixel <= "000000";
      when 19009 => pixel <= "000000";
      when 19010 => pixel <= "000000";
      when 19011 => pixel <= "000000";
      when 19012 => pixel <= "000000";
      when 19013 => pixel <= "000000";
      when 19014 => pixel <= "000000";
      when 19015 => pixel <= "000000";
      when 19016 => pixel <= "000000";
      when 19017 => pixel <= "000000";
      when 19018 => pixel <= "000000";
      when 19019 => pixel <= "000000";
      when 19020 => pixel <= "000000";
      when 19021 => pixel <= "000000";
      when 19022 => pixel <= "000000";
      when 19023 => pixel <= "000000";
      when 19024 => pixel <= "000000";
      when 19025 => pixel <= "000000";
      when 19026 => pixel <= "000000";
      when 19027 => pixel <= "000000";
      when 19028 => pixel <= "000000";
      when 19029 => pixel <= "000000";
      when 19030 => pixel <= "000000";
      when 19031 => pixel <= "000000";
      when 19032 => pixel <= "000000";
      when 19033 => pixel <= "000000";
      when 19034 => pixel <= "000000";
      when 19035 => pixel <= "000000";
      when 19036 => pixel <= "000000";
      when 19037 => pixel <= "000000";
      when 19038 => pixel <= "000000";
      when 19039 => pixel <= "000000";
      when 19040 => pixel <= "000000";
      when 19041 => pixel <= "000000";
      when 19042 => pixel <= "000000";
      when 19043 => pixel <= "000000";
      when 19044 => pixel <= "000000";
      when 19045 => pixel <= "000000";
      when 19046 => pixel <= "000000";
      when 19047 => pixel <= "000000";
      when 19048 => pixel <= "000000";
      when 19049 => pixel <= "000000";
      when 19050 => pixel <= "000000";
      when 19051 => pixel <= "000000";
      when 19052 => pixel <= "000000";
      when 19053 => pixel <= "000000";
      when 19054 => pixel <= "000000";
      when 19055 => pixel <= "000000";
      when 19056 => pixel <= "000000";
      when 19057 => pixel <= "000000";
      when 19058 => pixel <= "000000";
      when 19059 => pixel <= "000000";
      when 19060 => pixel <= "000000";
      when 19061 => pixel <= "000000";
      when 19062 => pixel <= "000000";
      when 19063 => pixel <= "000000";
      when 19064 => pixel <= "000000";
      when 19065 => pixel <= "000000";
      when 19066 => pixel <= "000000";
      when 19067 => pixel <= "000000";
      when 19068 => pixel <= "000000";
      when 19069 => pixel <= "000000";
      when 19070 => pixel <= "000000";
      when 19071 => pixel <= "000000";
      when 19072 => pixel <= "000000";
      when 19073 => pixel <= "000000";
      when 19074 => pixel <= "000000";
      when 19075 => pixel <= "000000";
      when 19076 => pixel <= "000000";
      when 19077 => pixel <= "000000";
      when 19078 => pixel <= "000000";
      when 19079 => pixel <= "000000";
      when 19080 => pixel <= "000000";
      when 19081 => pixel <= "000000";
      when 19082 => pixel <= "000000";
      when 19083 => pixel <= "000000";
      when 19084 => pixel <= "000000";
      when 19085 => pixel <= "000000";
      when 19086 => pixel <= "000000";
      when 19087 => pixel <= "000000";
      when 19088 => pixel <= "000000";
      when 19089 => pixel <= "000000";
      when 19090 => pixel <= "000000";
      when 19091 => pixel <= "000000";
      when 19092 => pixel <= "000000";
      when 19093 => pixel <= "000000";
      when 19094 => pixel <= "000000";
      when 19095 => pixel <= "000000";
      when 19096 => pixel <= "000000";
      when 19097 => pixel <= "000000";
      when 19098 => pixel <= "000000";
      when 19099 => pixel <= "000000";
      when 19100 => pixel <= "000000";
      when 19101 => pixel <= "000000";
      when 19102 => pixel <= "000000";
      when 19103 => pixel <= "000000";
      when 19104 => pixel <= "000000";
      when 19105 => pixel <= "000000";
      when 19106 => pixel <= "000000";
      when 19107 => pixel <= "000000";
      when 19108 => pixel <= "000000";
      when 19109 => pixel <= "000000";
      when 19110 => pixel <= "000000";
      when 19111 => pixel <= "000000";
      when 19112 => pixel <= "000000";
      when 19113 => pixel <= "000000";
      when 19114 => pixel <= "000000";
      when 19115 => pixel <= "000000";
      when 19116 => pixel <= "000000";
      when 19117 => pixel <= "000000";
      when 19118 => pixel <= "000000";
      when 19119 => pixel <= "000000";
      when 19120 => pixel <= "000000";
      when 19121 => pixel <= "000000";
      when 19122 => pixel <= "000000";
      when 19123 => pixel <= "000000";
      when 19124 => pixel <= "000000";
      when 19125 => pixel <= "000000";
      when 19126 => pixel <= "000000";
      when 19127 => pixel <= "000000";
      when 19128 => pixel <= "000000";
      when 19129 => pixel <= "000000";
      when 19130 => pixel <= "000000";
      when 19131 => pixel <= "000000";
      when 19132 => pixel <= "000000";
      when 19133 => pixel <= "000000";
      when 19134 => pixel <= "000000";
      when 19135 => pixel <= "000000";
      when 19136 => pixel <= "000000";
      when 19137 => pixel <= "000000";
      when 19138 => pixel <= "000000";
      when 19139 => pixel <= "000000";
      when 19140 => pixel <= "000000";
      when 19141 => pixel <= "000000";
      when 19142 => pixel <= "000000";
      when 19143 => pixel <= "000000";
      when 19144 => pixel <= "000000";
      when 19145 => pixel <= "000000";
      when 19146 => pixel <= "000000";
      when 19147 => pixel <= "000000";
      when 19148 => pixel <= "000000";
      when 19149 => pixel <= "000000";
      when 19150 => pixel <= "000000";
      when 19151 => pixel <= "000000";
      when 19152 => pixel <= "000000";
      when 19153 => pixel <= "000000";
      when 19154 => pixel <= "000000";
      when 19155 => pixel <= "000000";
      when 19156 => pixel <= "000000";
      when 19157 => pixel <= "000000";
      when 19158 => pixel <= "000000";
      when 19159 => pixel <= "000000";
      when 19160 => pixel <= "000000";
      when 19161 => pixel <= "000000";
      when 19162 => pixel <= "000000";
      when 19163 => pixel <= "000000";
      when 19164 => pixel <= "000000";
      when 19165 => pixel <= "000000";
      when 19166 => pixel <= "000000";
      when 19167 => pixel <= "000000";
      when 19168 => pixel <= "000000";
      when 19169 => pixel <= "000000";
      when 19170 => pixel <= "000000";
      when 19171 => pixel <= "000000";
      when 19172 => pixel <= "000000";
      when 19173 => pixel <= "000000";
      when 19174 => pixel <= "000000";
      when 19175 => pixel <= "000000";
      when 19176 => pixel <= "000000";
      when 19177 => pixel <= "000000";
      when 19178 => pixel <= "000000";
      when 19179 => pixel <= "000000";
      when 19180 => pixel <= "000000";
      when 19181 => pixel <= "000000";
      when 19182 => pixel <= "000000";
      when 19183 => pixel <= "000000";
      when 19184 => pixel <= "000000";
      when 19185 => pixel <= "000000";
      when 19186 => pixel <= "000000";
      when 19187 => pixel <= "000000";
      when 19188 => pixel <= "000000";
      when 19189 => pixel <= "000000";
      when 19190 => pixel <= "000000";
      when 19191 => pixel <= "000000";
      when 19192 => pixel <= "000000";
      when 19193 => pixel <= "000000";
      when 19194 => pixel <= "000000";
      when 19195 => pixel <= "000000";
      when 19196 => pixel <= "000000";
      when 19197 => pixel <= "000000";
      when 19198 => pixel <= "000000";
      when 19199 => pixel <= "000000";
      when others => pixel <= (others => '0');
    end case;
  end process;
end;

