library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity numbers_rom is
  port (
    x     : in  std_logic_vector(7 downto 0);
    y     : in  std_logic_vector(3 downto 0);
    pixel : out std_logic_vector(5 downto 0)
  );
end entity;

architecture synth of numbers_rom is
  signal addr : unsigned(11 downto 0);
begin
  addr <= (unsigned(y) * 8d"160") + unsigned(x);
  process(addr)
  begin
    case addr is
      when 0 => pixel <= "111111";
      when 1 => pixel <= "111111";
      when 2 => pixel <= "111111";
      when 3 => pixel <= "111111";
      when 4 => pixel <= "111111";
      when 5 => pixel <= "111111";
      when 6 => pixel <= "111111";
      when 7 => pixel <= "111111";
      when 8 => pixel <= "111111";
      when 9 => pixel <= "111111";
      when 10 => pixel <= "111111";
      when 11 => pixel <= "111111";
      when 12 => pixel <= "111111";
      when 13 => pixel <= "111111";
      when 14 => pixel <= "111111";
      when 15 => pixel <= "111111";
      when 16 => pixel <= "111111";
      when 17 => pixel <= "111111";
      when 18 => pixel <= "111111";
      when 19 => pixel <= "111111";
      when 20 => pixel <= "111111";
      when 21 => pixel <= "111111";
      when 22 => pixel <= "111111";
      when 23 => pixel <= "111111";
      when 24 => pixel <= "111111";
      when 25 => pixel <= "111111";
      when 26 => pixel <= "111111";
      when 27 => pixel <= "111111";
      when 28 => pixel <= "111111";
      when 29 => pixel <= "111111";
      when 30 => pixel <= "111111";
      when 31 => pixel <= "111111";
      when 32 => pixel <= "111111";
      when 33 => pixel <= "111111";
      when 34 => pixel <= "111111";
      when 35 => pixel <= "111111";
      when 36 => pixel <= "111111";
      when 37 => pixel <= "111111";
      when 38 => pixel <= "111111";
      when 39 => pixel <= "111111";
      when 40 => pixel <= "111111";
      when 41 => pixel <= "111111";
      when 42 => pixel <= "111111";
      when 43 => pixel <= "111111";
      when 44 => pixel <= "111111";
      when 45 => pixel <= "111111";
      when 46 => pixel <= "111111";
      when 47 => pixel <= "111111";
      when 48 => pixel <= "111111";
      when 49 => pixel <= "111111";
      when 50 => pixel <= "111111";
      when 51 => pixel <= "111111";
      when 52 => pixel <= "111111";
      when 53 => pixel <= "111111";
      when 54 => pixel <= "111111";
      when 55 => pixel <= "111111";
      when 56 => pixel <= "111111";
      when 57 => pixel <= "111111";
      when 58 => pixel <= "111111";
      when 59 => pixel <= "111111";
      when 60 => pixel <= "111111";
      when 61 => pixel <= "111111";
      when 62 => pixel <= "111111";
      when 63 => pixel <= "111111";
      when 64 => pixel <= "111111";
      when 65 => pixel <= "111111";
      when 66 => pixel <= "111111";
      when 67 => pixel <= "111111";
      when 68 => pixel <= "111111";
      when 69 => pixel <= "111111";
      when 70 => pixel <= "111111";
      when 71 => pixel <= "111111";
      when 72 => pixel <= "111111";
      when 73 => pixel <= "111111";
      when 74 => pixel <= "111111";
      when 75 => pixel <= "111111";
      when 76 => pixel <= "111111";
      when 77 => pixel <= "111111";
      when 78 => pixel <= "111111";
      when 79 => pixel <= "111111";
      when 80 => pixel <= "111111";
      when 81 => pixel <= "111111";
      when 82 => pixel <= "111111";
      when 83 => pixel <= "111111";
      when 84 => pixel <= "111111";
      when 85 => pixel <= "111111";
      when 86 => pixel <= "111111";
      when 87 => pixel <= "111111";
      when 88 => pixel <= "111111";
      when 89 => pixel <= "111111";
      when 90 => pixel <= "111111";
      when 91 => pixel <= "111111";
      when 92 => pixel <= "111111";
      when 93 => pixel <= "111111";
      when 94 => pixel <= "111111";
      when 95 => pixel <= "111111";
      when 96 => pixel <= "111111";
      when 97 => pixel <= "111111";
      when 98 => pixel <= "111111";
      when 99 => pixel <= "111111";
      when 100 => pixel <= "111111";
      when 101 => pixel <= "111111";
      when 102 => pixel <= "111111";
      when 103 => pixel <= "111111";
      when 104 => pixel <= "111111";
      when 105 => pixel <= "111111";
      when 106 => pixel <= "111111";
      when 107 => pixel <= "111111";
      when 108 => pixel <= "111111";
      when 109 => pixel <= "111111";
      when 110 => pixel <= "111111";
      when 111 => pixel <= "111111";
      when 112 => pixel <= "111111";
      when 113 => pixel <= "111111";
      when 114 => pixel <= "111111";
      when 115 => pixel <= "111111";
      when 116 => pixel <= "111111";
      when 117 => pixel <= "111111";
      when 118 => pixel <= "111111";
      when 119 => pixel <= "111111";
      when 120 => pixel <= "111111";
      when 121 => pixel <= "111111";
      when 122 => pixel <= "111111";
      when 123 => pixel <= "111111";
      when 124 => pixel <= "111111";
      when 125 => pixel <= "111111";
      when 126 => pixel <= "111111";
      when 127 => pixel <= "111111";
      when 128 => pixel <= "111111";
      when 129 => pixel <= "111111";
      when 130 => pixel <= "111111";
      when 131 => pixel <= "111111";
      when 132 => pixel <= "111111";
      when 133 => pixel <= "111111";
      when 134 => pixel <= "111111";
      when 135 => pixel <= "111111";
      when 136 => pixel <= "111111";
      when 137 => pixel <= "111111";
      when 138 => pixel <= "111111";
      when 139 => pixel <= "111111";
      when 140 => pixel <= "111111";
      when 141 => pixel <= "111111";
      when 142 => pixel <= "111111";
      when 143 => pixel <= "111111";
      when 144 => pixel <= "111111";
      when 145 => pixel <= "111111";
      when 146 => pixel <= "111111";
      when 147 => pixel <= "111111";
      when 148 => pixel <= "111111";
      when 149 => pixel <= "111111";
      when 150 => pixel <= "111111";
      when 151 => pixel <= "111111";
      when 152 => pixel <= "111111";
      when 153 => pixel <= "111111";
      when 154 => pixel <= "111111";
      when 155 => pixel <= "111111";
      when 156 => pixel <= "111111";
      when 157 => pixel <= "111111";
      when 158 => pixel <= "111111";
      when 159 => pixel <= "111111";
      when 160 => pixel <= "111111";
      when 161 => pixel <= "111111";
      when 162 => pixel <= "111111";
      when 163 => pixel <= "111111";
      when 164 => pixel <= "111111";
      when 165 => pixel <= "111111";
      when 166 => pixel <= "111111";
      when 167 => pixel <= "111111";
      when 168 => pixel <= "111111";
      when 169 => pixel <= "111111";
      when 170 => pixel <= "111111";
      when 171 => pixel <= "111111";
      when 172 => pixel <= "111111";
      when 173 => pixel <= "111111";
      when 174 => pixel <= "111111";
      when 175 => pixel <= "111111";
      when 176 => pixel <= "111111";
      when 177 => pixel <= "111111";
      when 178 => pixel <= "111111";
      when 179 => pixel <= "111111";
      when 180 => pixel <= "111111";
      when 181 => pixel <= "111111";
      when 182 => pixel <= "111111";
      when 183 => pixel <= "111111";
      when 184 => pixel <= "111111";
      when 185 => pixel <= "111111";
      when 186 => pixel <= "111111";
      when 187 => pixel <= "111111";
      when 188 => pixel <= "111111";
      when 189 => pixel <= "111111";
      when 190 => pixel <= "111111";
      when 191 => pixel <= "111111";
      when 192 => pixel <= "111111";
      when 193 => pixel <= "111111";
      when 194 => pixel <= "111111";
      when 195 => pixel <= "111111";
      when 196 => pixel <= "111111";
      when 197 => pixel <= "111111";
      when 198 => pixel <= "111111";
      when 199 => pixel <= "111111";
      when 200 => pixel <= "111111";
      when 201 => pixel <= "111111";
      when 202 => pixel <= "111111";
      when 203 => pixel <= "111111";
      when 204 => pixel <= "111111";
      when 205 => pixel <= "111111";
      when 206 => pixel <= "111111";
      when 207 => pixel <= "111111";
      when 208 => pixel <= "111111";
      when 209 => pixel <= "111111";
      when 210 => pixel <= "111111";
      when 211 => pixel <= "111111";
      when 212 => pixel <= "111111";
      when 213 => pixel <= "111111";
      when 214 => pixel <= "111111";
      when 215 => pixel <= "111111";
      when 216 => pixel <= "111111";
      when 217 => pixel <= "111111";
      when 218 => pixel <= "111111";
      when 219 => pixel <= "111111";
      when 220 => pixel <= "111111";
      when 221 => pixel <= "111111";
      when 222 => pixel <= "111111";
      when 223 => pixel <= "111111";
      when 224 => pixel <= "111111";
      when 225 => pixel <= "111111";
      when 226 => pixel <= "111111";
      when 227 => pixel <= "111111";
      when 228 => pixel <= "111111";
      when 229 => pixel <= "111111";
      when 230 => pixel <= "111111";
      when 231 => pixel <= "111111";
      when 232 => pixel <= "111111";
      when 233 => pixel <= "111111";
      when 234 => pixel <= "111111";
      when 235 => pixel <= "111111";
      when 236 => pixel <= "111111";
      when 237 => pixel <= "111111";
      when 238 => pixel <= "111111";
      when 239 => pixel <= "111111";
      when 240 => pixel <= "111111";
      when 241 => pixel <= "111111";
      when 242 => pixel <= "111111";
      when 243 => pixel <= "111111";
      when 244 => pixel <= "111111";
      when 245 => pixel <= "111111";
      when 246 => pixel <= "111111";
      when 247 => pixel <= "111111";
      when 248 => pixel <= "111111";
      when 249 => pixel <= "111111";
      when 250 => pixel <= "111111";
      when 251 => pixel <= "111111";
      when 252 => pixel <= "111111";
      when 253 => pixel <= "111111";
      when 254 => pixel <= "111111";
      when 255 => pixel <= "111111";
      when 256 => pixel <= "111111";
      when 257 => pixel <= "111111";
      when 258 => pixel <= "111111";
      when 259 => pixel <= "111111";
      when 260 => pixel <= "111111";
      when 261 => pixel <= "111111";
      when 262 => pixel <= "111111";
      when 263 => pixel <= "111111";
      when 264 => pixel <= "111111";
      when 265 => pixel <= "111111";
      when 266 => pixel <= "111111";
      when 267 => pixel <= "111111";
      when 268 => pixel <= "111111";
      when 269 => pixel <= "111111";
      when 270 => pixel <= "111111";
      when 271 => pixel <= "111111";
      when 272 => pixel <= "111111";
      when 273 => pixel <= "111111";
      when 274 => pixel <= "111111";
      when 275 => pixel <= "111111";
      when 276 => pixel <= "111111";
      when 277 => pixel <= "111111";
      when 278 => pixel <= "111111";
      when 279 => pixel <= "111111";
      when 280 => pixel <= "111111";
      when 281 => pixel <= "111111";
      when 282 => pixel <= "111111";
      when 283 => pixel <= "111111";
      when 284 => pixel <= "111111";
      when 285 => pixel <= "111111";
      when 286 => pixel <= "111111";
      when 287 => pixel <= "111111";
      when 288 => pixel <= "111111";
      when 289 => pixel <= "111111";
      when 290 => pixel <= "111111";
      when 291 => pixel <= "111111";
      when 292 => pixel <= "111111";
      when 293 => pixel <= "111111";
      when 294 => pixel <= "111111";
      when 295 => pixel <= "111111";
      when 296 => pixel <= "111111";
      when 297 => pixel <= "111111";
      when 298 => pixel <= "111111";
      when 299 => pixel <= "111111";
      when 300 => pixel <= "111111";
      when 301 => pixel <= "111111";
      when 302 => pixel <= "111111";
      when 303 => pixel <= "111111";
      when 304 => pixel <= "111111";
      when 305 => pixel <= "111111";
      when 306 => pixel <= "111111";
      when 307 => pixel <= "111111";
      when 308 => pixel <= "111111";
      when 309 => pixel <= "111111";
      when 310 => pixel <= "111111";
      when 311 => pixel <= "111111";
      when 312 => pixel <= "111111";
      when 313 => pixel <= "111111";
      when 314 => pixel <= "111111";
      when 315 => pixel <= "111111";
      when 316 => pixel <= "111111";
      when 317 => pixel <= "111111";
      when 318 => pixel <= "111111";
      when 319 => pixel <= "111111";
      when 320 => pixel <= "111111";
      when 321 => pixel <= "111111";
      when 322 => pixel <= "111111";
      when 323 => pixel <= "111111";
      when 324 => pixel <= "111111";
      when 325 => pixel <= "111111";
      when 326 => pixel <= "111111";
      when 327 => pixel <= "111111";
      when 328 => pixel <= "111111";
      when 329 => pixel <= "111111";
      when 330 => pixel <= "111111";
      when 331 => pixel <= "111111";
      when 332 => pixel <= "111111";
      when 333 => pixel <= "111111";
      when 334 => pixel <= "111111";
      when 335 => pixel <= "111111";
      when 336 => pixel <= "111111";
      when 337 => pixel <= "111111";
      when 338 => pixel <= "111111";
      when 339 => pixel <= "111111";
      when 340 => pixel <= "111111";
      when 341 => pixel <= "111111";
      when 342 => pixel <= "111111";
      when 343 => pixel <= "111111";
      when 344 => pixel <= "111111";
      when 345 => pixel <= "111111";
      when 346 => pixel <= "111111";
      when 347 => pixel <= "111111";
      when 348 => pixel <= "111111";
      when 349 => pixel <= "111111";
      when 350 => pixel <= "111111";
      when 351 => pixel <= "111111";
      when 352 => pixel <= "111111";
      when 353 => pixel <= "111111";
      when 354 => pixel <= "111111";
      when 355 => pixel <= "111111";
      when 356 => pixel <= "111111";
      when 357 => pixel <= "111111";
      when 358 => pixel <= "111111";
      when 359 => pixel <= "111111";
      when 360 => pixel <= "111111";
      when 361 => pixel <= "111111";
      when 362 => pixel <= "111111";
      when 363 => pixel <= "111111";
      when 364 => pixel <= "111111";
      when 365 => pixel <= "111111";
      when 366 => pixel <= "111111";
      when 367 => pixel <= "111111";
      when 368 => pixel <= "111111";
      when 369 => pixel <= "111111";
      when 370 => pixel <= "111111";
      when 371 => pixel <= "111111";
      when 372 => pixel <= "111111";
      when 373 => pixel <= "111111";
      when 374 => pixel <= "111111";
      when 375 => pixel <= "111111";
      when 376 => pixel <= "111111";
      when 377 => pixel <= "111111";
      when 378 => pixel <= "111111";
      when 379 => pixel <= "111111";
      when 380 => pixel <= "111111";
      when 381 => pixel <= "111111";
      when 382 => pixel <= "111111";
      when 383 => pixel <= "111111";
      when 384 => pixel <= "111111";
      when 385 => pixel <= "111111";
      when 386 => pixel <= "111111";
      when 387 => pixel <= "111111";
      when 388 => pixel <= "111111";
      when 389 => pixel <= "111111";
      when 390 => pixel <= "111111";
      when 391 => pixel <= "111111";
      when 392 => pixel <= "111111";
      when 393 => pixel <= "111111";
      when 394 => pixel <= "111111";
      when 395 => pixel <= "111111";
      when 396 => pixel <= "111111";
      when 397 => pixel <= "111111";
      when 398 => pixel <= "111111";
      when 399 => pixel <= "111111";
      when 400 => pixel <= "111111";
      when 401 => pixel <= "111111";
      when 402 => pixel <= "111111";
      when 403 => pixel <= "111111";
      when 404 => pixel <= "111111";
      when 405 => pixel <= "111111";
      when 406 => pixel <= "111111";
      when 407 => pixel <= "111111";
      when 408 => pixel <= "111111";
      when 409 => pixel <= "111111";
      when 410 => pixel <= "111111";
      when 411 => pixel <= "111111";
      when 412 => pixel <= "111111";
      when 413 => pixel <= "111111";
      when 414 => pixel <= "111111";
      when 415 => pixel <= "111111";
      when 416 => pixel <= "111111";
      when 417 => pixel <= "111111";
      when 418 => pixel <= "111111";
      when 419 => pixel <= "111111";
      when 420 => pixel <= "111111";
      when 421 => pixel <= "111111";
      when 422 => pixel <= "111111";
      when 423 => pixel <= "111111";
      when 424 => pixel <= "111111";
      when 425 => pixel <= "111111";
      when 426 => pixel <= "111111";
      when 427 => pixel <= "111111";
      when 428 => pixel <= "111111";
      when 429 => pixel <= "111111";
      when 430 => pixel <= "111111";
      when 431 => pixel <= "111111";
      when 432 => pixel <= "111111";
      when 433 => pixel <= "111111";
      when 434 => pixel <= "111111";
      when 435 => pixel <= "111111";
      when 436 => pixel <= "111111";
      when 437 => pixel <= "111111";
      when 438 => pixel <= "111111";
      when 439 => pixel <= "111111";
      when 440 => pixel <= "111111";
      when 441 => pixel <= "111111";
      when 442 => pixel <= "111111";
      when 443 => pixel <= "111111";
      when 444 => pixel <= "111111";
      when 445 => pixel <= "111111";
      when 446 => pixel <= "111111";
      when 447 => pixel <= "111111";
      when 448 => pixel <= "111111";
      when 449 => pixel <= "111111";
      when 450 => pixel <= "111111";
      when 451 => pixel <= "111111";
      when 452 => pixel <= "111111";
      when 453 => pixel <= "111111";
      when 454 => pixel <= "111111";
      when 455 => pixel <= "111111";
      when 456 => pixel <= "111111";
      when 457 => pixel <= "111111";
      when 458 => pixel <= "111111";
      when 459 => pixel <= "111111";
      when 460 => pixel <= "111111";
      when 461 => pixel <= "111111";
      when 462 => pixel <= "111111";
      when 463 => pixel <= "111111";
      when 464 => pixel <= "111111";
      when 465 => pixel <= "111111";
      when 466 => pixel <= "111111";
      when 467 => pixel <= "111111";
      when 468 => pixel <= "111111";
      when 469 => pixel <= "111111";
      when 470 => pixel <= "111111";
      when 471 => pixel <= "111111";
      when 472 => pixel <= "111111";
      when 473 => pixel <= "111111";
      when 474 => pixel <= "111111";
      when 475 => pixel <= "111111";
      when 476 => pixel <= "111111";
      when 477 => pixel <= "111111";
      when 478 => pixel <= "111111";
      when 479 => pixel <= "111111";
      when 480 => pixel <= "111111";
      when 481 => pixel <= "111111";
      when 482 => pixel <= "111111";
      when 483 => pixel <= "111111";
      when 484 => pixel <= "111111";
      when 485 => pixel <= "111111";
      when 486 => pixel <= "000000";
      when 487 => pixel <= "000000";
      when 488 => pixel <= "000000";
      when 489 => pixel <= "111111";
      when 490 => pixel <= "111111";
      when 491 => pixel <= "111111";
      when 492 => pixel <= "111111";
      when 493 => pixel <= "111111";
      when 494 => pixel <= "111111";
      when 495 => pixel <= "111111";
      when 496 => pixel <= "111111";
      when 497 => pixel <= "111111";
      when 498 => pixel <= "111111";
      when 499 => pixel <= "111111";
      when 500 => pixel <= "111111";
      when 501 => pixel <= "111111";
      when 502 => pixel <= "111111";
      when 503 => pixel <= "000000";
      when 504 => pixel <= "000000";
      when 505 => pixel <= "111111";
      when 506 => pixel <= "111111";
      when 507 => pixel <= "111111";
      when 508 => pixel <= "111111";
      when 509 => pixel <= "111111";
      when 510 => pixel <= "111111";
      when 511 => pixel <= "111111";
      when 512 => pixel <= "111111";
      when 513 => pixel <= "111111";
      when 514 => pixel <= "111111";
      when 515 => pixel <= "111111";
      when 516 => pixel <= "111111";
      when 517 => pixel <= "000000";
      when 518 => pixel <= "000000";
      when 519 => pixel <= "000000";
      when 520 => pixel <= "000000";
      when 521 => pixel <= "000000";
      when 522 => pixel <= "111111";
      when 523 => pixel <= "111111";
      when 524 => pixel <= "111111";
      when 525 => pixel <= "111111";
      when 526 => pixel <= "111111";
      when 527 => pixel <= "111111";
      when 528 => pixel <= "111111";
      when 529 => pixel <= "111111";
      when 530 => pixel <= "111111";
      when 531 => pixel <= "111111";
      when 532 => pixel <= "111111";
      when 533 => pixel <= "000000";
      when 534 => pixel <= "000000";
      when 535 => pixel <= "000000";
      when 536 => pixel <= "000000";
      when 537 => pixel <= "000000";
      when 538 => pixel <= "111111";
      when 539 => pixel <= "111111";
      when 540 => pixel <= "111111";
      when 541 => pixel <= "111111";
      when 542 => pixel <= "111111";
      when 543 => pixel <= "111111";
      when 544 => pixel <= "111111";
      when 545 => pixel <= "111111";
      when 546 => pixel <= "111111";
      when 547 => pixel <= "111111";
      when 548 => pixel <= "111111";
      when 549 => pixel <= "111111";
      when 550 => pixel <= "111111";
      when 551 => pixel <= "111111";
      when 552 => pixel <= "000000";
      when 553 => pixel <= "000000";
      when 554 => pixel <= "111111";
      when 555 => pixel <= "111111";
      when 556 => pixel <= "111111";
      when 557 => pixel <= "111111";
      when 558 => pixel <= "111111";
      when 559 => pixel <= "111111";
      when 560 => pixel <= "111111";
      when 561 => pixel <= "111111";
      when 562 => pixel <= "111111";
      when 563 => pixel <= "111111";
      when 564 => pixel <= "000000";
      when 565 => pixel <= "000000";
      when 566 => pixel <= "000000";
      when 567 => pixel <= "000000";
      when 568 => pixel <= "000000";
      when 569 => pixel <= "000000";
      when 570 => pixel <= "000000";
      when 571 => pixel <= "111111";
      when 572 => pixel <= "111111";
      when 573 => pixel <= "111111";
      when 574 => pixel <= "111111";
      when 575 => pixel <= "111111";
      when 576 => pixel <= "111111";
      when 577 => pixel <= "111111";
      when 578 => pixel <= "111111";
      when 579 => pixel <= "111111";
      when 580 => pixel <= "111111";
      when 581 => pixel <= "111111";
      when 582 => pixel <= "000000";
      when 583 => pixel <= "000000";
      when 584 => pixel <= "000000";
      when 585 => pixel <= "111111";
      when 586 => pixel <= "111111";
      when 587 => pixel <= "111111";
      when 588 => pixel <= "111111";
      when 589 => pixel <= "111111";
      when 590 => pixel <= "111111";
      when 591 => pixel <= "111111";
      when 592 => pixel <= "111111";
      when 593 => pixel <= "111111";
      when 594 => pixel <= "111111";
      when 595 => pixel <= "111111";
      when 596 => pixel <= "000000";
      when 597 => pixel <= "000000";
      when 598 => pixel <= "000000";
      when 599 => pixel <= "000000";
      when 600 => pixel <= "000000";
      when 601 => pixel <= "000000";
      when 602 => pixel <= "000000";
      when 603 => pixel <= "111111";
      when 604 => pixel <= "111111";
      when 605 => pixel <= "111111";
      when 606 => pixel <= "111111";
      when 607 => pixel <= "111111";
      when 608 => pixel <= "111111";
      when 609 => pixel <= "111111";
      when 610 => pixel <= "111111";
      when 611 => pixel <= "111111";
      when 612 => pixel <= "111111";
      when 613 => pixel <= "000000";
      when 614 => pixel <= "000000";
      when 615 => pixel <= "000000";
      when 616 => pixel <= "000000";
      when 617 => pixel <= "000000";
      when 618 => pixel <= "111111";
      when 619 => pixel <= "111111";
      when 620 => pixel <= "111111";
      when 621 => pixel <= "111111";
      when 622 => pixel <= "111111";
      when 623 => pixel <= "111111";
      when 624 => pixel <= "111111";
      when 625 => pixel <= "111111";
      when 626 => pixel <= "111111";
      when 627 => pixel <= "111111";
      when 628 => pixel <= "111111";
      when 629 => pixel <= "000000";
      when 630 => pixel <= "000000";
      when 631 => pixel <= "000000";
      when 632 => pixel <= "000000";
      when 633 => pixel <= "000000";
      when 634 => pixel <= "111111";
      when 635 => pixel <= "111111";
      when 636 => pixel <= "111111";
      when 637 => pixel <= "111111";
      when 638 => pixel <= "111111";
      when 639 => pixel <= "111111";
      when 640 => pixel <= "111111";
      when 641 => pixel <= "111111";
      when 642 => pixel <= "111111";
      when 643 => pixel <= "111111";
      when 644 => pixel <= "111111";
      when 645 => pixel <= "000000";
      when 646 => pixel <= "000000";
      when 647 => pixel <= "111111";
      when 648 => pixel <= "000000";
      when 649 => pixel <= "000000";
      when 650 => pixel <= "111111";
      when 651 => pixel <= "111111";
      when 652 => pixel <= "111111";
      when 653 => pixel <= "111111";
      when 654 => pixel <= "111111";
      when 655 => pixel <= "111111";
      when 656 => pixel <= "111111";
      when 657 => pixel <= "111111";
      when 658 => pixel <= "111111";
      when 659 => pixel <= "111111";
      when 660 => pixel <= "111111";
      when 661 => pixel <= "111111";
      when 662 => pixel <= "000000";
      when 663 => pixel <= "000000";
      when 664 => pixel <= "000000";
      when 665 => pixel <= "111111";
      when 666 => pixel <= "111111";
      when 667 => pixel <= "111111";
      when 668 => pixel <= "111111";
      when 669 => pixel <= "111111";
      when 670 => pixel <= "111111";
      when 671 => pixel <= "111111";
      when 672 => pixel <= "111111";
      when 673 => pixel <= "111111";
      when 674 => pixel <= "111111";
      when 675 => pixel <= "111111";
      when 676 => pixel <= "000000";
      when 677 => pixel <= "000000";
      when 678 => pixel <= "111111";
      when 679 => pixel <= "111111";
      when 680 => pixel <= "111111";
      when 681 => pixel <= "000000";
      when 682 => pixel <= "000000";
      when 683 => pixel <= "111111";
      when 684 => pixel <= "111111";
      when 685 => pixel <= "111111";
      when 686 => pixel <= "111111";
      when 687 => pixel <= "111111";
      when 688 => pixel <= "111111";
      when 689 => pixel <= "111111";
      when 690 => pixel <= "111111";
      when 691 => pixel <= "111111";
      when 692 => pixel <= "000000";
      when 693 => pixel <= "000000";
      when 694 => pixel <= "111111";
      when 695 => pixel <= "111111";
      when 696 => pixel <= "111111";
      when 697 => pixel <= "000000";
      when 698 => pixel <= "000000";
      when 699 => pixel <= "111111";
      when 700 => pixel <= "111111";
      when 701 => pixel <= "111111";
      when 702 => pixel <= "111111";
      when 703 => pixel <= "111111";
      when 704 => pixel <= "111111";
      when 705 => pixel <= "111111";
      when 706 => pixel <= "111111";
      when 707 => pixel <= "111111";
      when 708 => pixel <= "111111";
      when 709 => pixel <= "111111";
      when 710 => pixel <= "111111";
      when 711 => pixel <= "000000";
      when 712 => pixel <= "000000";
      when 713 => pixel <= "000000";
      when 714 => pixel <= "111111";
      when 715 => pixel <= "111111";
      when 716 => pixel <= "111111";
      when 717 => pixel <= "111111";
      when 718 => pixel <= "111111";
      when 719 => pixel <= "111111";
      when 720 => pixel <= "111111";
      when 721 => pixel <= "111111";
      when 722 => pixel <= "111111";
      when 723 => pixel <= "111111";
      when 724 => pixel <= "000000";
      when 725 => pixel <= "000000";
      when 726 => pixel <= "111111";
      when 727 => pixel <= "111111";
      when 728 => pixel <= "111111";
      when 729 => pixel <= "111111";
      when 730 => pixel <= "111111";
      when 731 => pixel <= "111111";
      when 732 => pixel <= "111111";
      when 733 => pixel <= "111111";
      when 734 => pixel <= "111111";
      when 735 => pixel <= "111111";
      when 736 => pixel <= "111111";
      when 737 => pixel <= "111111";
      when 738 => pixel <= "111111";
      when 739 => pixel <= "111111";
      when 740 => pixel <= "111111";
      when 741 => pixel <= "000000";
      when 742 => pixel <= "000000";
      when 743 => pixel <= "111111";
      when 744 => pixel <= "111111";
      when 745 => pixel <= "111111";
      when 746 => pixel <= "111111";
      when 747 => pixel <= "111111";
      when 748 => pixel <= "111111";
      when 749 => pixel <= "111111";
      when 750 => pixel <= "111111";
      when 751 => pixel <= "111111";
      when 752 => pixel <= "111111";
      when 753 => pixel <= "111111";
      when 754 => pixel <= "111111";
      when 755 => pixel <= "111111";
      when 756 => pixel <= "000000";
      when 757 => pixel <= "000000";
      when 758 => pixel <= "111111";
      when 759 => pixel <= "111111";
      when 760 => pixel <= "111111";
      when 761 => pixel <= "000000";
      when 762 => pixel <= "000000";
      when 763 => pixel <= "111111";
      when 764 => pixel <= "111111";
      when 765 => pixel <= "111111";
      when 766 => pixel <= "111111";
      when 767 => pixel <= "111111";
      when 768 => pixel <= "111111";
      when 769 => pixel <= "111111";
      when 770 => pixel <= "111111";
      when 771 => pixel <= "111111";
      when 772 => pixel <= "000000";
      when 773 => pixel <= "000000";
      when 774 => pixel <= "111111";
      when 775 => pixel <= "111111";
      when 776 => pixel <= "111111";
      when 777 => pixel <= "000000";
      when 778 => pixel <= "000000";
      when 779 => pixel <= "111111";
      when 780 => pixel <= "111111";
      when 781 => pixel <= "111111";
      when 782 => pixel <= "111111";
      when 783 => pixel <= "111111";
      when 784 => pixel <= "111111";
      when 785 => pixel <= "111111";
      when 786 => pixel <= "111111";
      when 787 => pixel <= "111111";
      when 788 => pixel <= "000000";
      when 789 => pixel <= "000000";
      when 790 => pixel <= "111111";
      when 791 => pixel <= "111111";
      when 792 => pixel <= "111111";
      when 793 => pixel <= "000000";
      when 794 => pixel <= "000000";
      when 795 => pixel <= "111111";
      when 796 => pixel <= "111111";
      when 797 => pixel <= "111111";
      when 798 => pixel <= "111111";
      when 799 => pixel <= "111111";
      when 800 => pixel <= "111111";
      when 801 => pixel <= "111111";
      when 802 => pixel <= "111111";
      when 803 => pixel <= "111111";
      when 804 => pixel <= "000000";
      when 805 => pixel <= "000000";
      when 806 => pixel <= "111111";
      when 807 => pixel <= "111111";
      when 808 => pixel <= "111111";
      when 809 => pixel <= "000000";
      when 810 => pixel <= "000000";
      when 811 => pixel <= "111111";
      when 812 => pixel <= "111111";
      when 813 => pixel <= "111111";
      when 814 => pixel <= "111111";
      when 815 => pixel <= "111111";
      when 816 => pixel <= "111111";
      when 817 => pixel <= "111111";
      when 818 => pixel <= "111111";
      when 819 => pixel <= "111111";
      when 820 => pixel <= "111111";
      when 821 => pixel <= "000000";
      when 822 => pixel <= "000000";
      when 823 => pixel <= "000000";
      when 824 => pixel <= "000000";
      when 825 => pixel <= "111111";
      when 826 => pixel <= "111111";
      when 827 => pixel <= "111111";
      when 828 => pixel <= "111111";
      when 829 => pixel <= "111111";
      when 830 => pixel <= "111111";
      when 831 => pixel <= "111111";
      when 832 => pixel <= "111111";
      when 833 => pixel <= "111111";
      when 834 => pixel <= "111111";
      when 835 => pixel <= "111111";
      when 836 => pixel <= "111111";
      when 837 => pixel <= "111111";
      when 838 => pixel <= "111111";
      when 839 => pixel <= "111111";
      when 840 => pixel <= "111111";
      when 841 => pixel <= "000000";
      when 842 => pixel <= "000000";
      when 843 => pixel <= "111111";
      when 844 => pixel <= "111111";
      when 845 => pixel <= "111111";
      when 846 => pixel <= "111111";
      when 847 => pixel <= "111111";
      when 848 => pixel <= "111111";
      when 849 => pixel <= "111111";
      when 850 => pixel <= "111111";
      when 851 => pixel <= "111111";
      when 852 => pixel <= "111111";
      when 853 => pixel <= "111111";
      when 854 => pixel <= "111111";
      when 855 => pixel <= "111111";
      when 856 => pixel <= "111111";
      when 857 => pixel <= "000000";
      when 858 => pixel <= "000000";
      when 859 => pixel <= "111111";
      when 860 => pixel <= "111111";
      when 861 => pixel <= "111111";
      when 862 => pixel <= "111111";
      when 863 => pixel <= "111111";
      when 864 => pixel <= "111111";
      when 865 => pixel <= "111111";
      when 866 => pixel <= "111111";
      when 867 => pixel <= "111111";
      when 868 => pixel <= "111111";
      when 869 => pixel <= "111111";
      when 870 => pixel <= "000000";
      when 871 => pixel <= "000000";
      when 872 => pixel <= "000000";
      when 873 => pixel <= "000000";
      when 874 => pixel <= "111111";
      when 875 => pixel <= "111111";
      when 876 => pixel <= "111111";
      when 877 => pixel <= "111111";
      when 878 => pixel <= "111111";
      when 879 => pixel <= "111111";
      when 880 => pixel <= "111111";
      when 881 => pixel <= "111111";
      when 882 => pixel <= "111111";
      when 883 => pixel <= "111111";
      when 884 => pixel <= "000000";
      when 885 => pixel <= "000000";
      when 886 => pixel <= "111111";
      when 887 => pixel <= "111111";
      when 888 => pixel <= "111111";
      when 889 => pixel <= "111111";
      when 890 => pixel <= "111111";
      when 891 => pixel <= "111111";
      when 892 => pixel <= "111111";
      when 893 => pixel <= "111111";
      when 894 => pixel <= "111111";
      when 895 => pixel <= "111111";
      when 896 => pixel <= "111111";
      when 897 => pixel <= "111111";
      when 898 => pixel <= "111111";
      when 899 => pixel <= "111111";
      when 900 => pixel <= "000000";
      when 901 => pixel <= "000000";
      when 902 => pixel <= "111111";
      when 903 => pixel <= "111111";
      when 904 => pixel <= "111111";
      when 905 => pixel <= "111111";
      when 906 => pixel <= "111111";
      when 907 => pixel <= "111111";
      when 908 => pixel <= "111111";
      when 909 => pixel <= "111111";
      when 910 => pixel <= "111111";
      when 911 => pixel <= "111111";
      when 912 => pixel <= "111111";
      when 913 => pixel <= "111111";
      when 914 => pixel <= "111111";
      when 915 => pixel <= "111111";
      when 916 => pixel <= "111111";
      when 917 => pixel <= "111111";
      when 918 => pixel <= "111111";
      when 919 => pixel <= "111111";
      when 920 => pixel <= "111111";
      when 921 => pixel <= "000000";
      when 922 => pixel <= "000000";
      when 923 => pixel <= "111111";
      when 924 => pixel <= "111111";
      when 925 => pixel <= "111111";
      when 926 => pixel <= "111111";
      when 927 => pixel <= "111111";
      when 928 => pixel <= "111111";
      when 929 => pixel <= "111111";
      when 930 => pixel <= "111111";
      when 931 => pixel <= "111111";
      when 932 => pixel <= "000000";
      when 933 => pixel <= "000000";
      when 934 => pixel <= "111111";
      when 935 => pixel <= "111111";
      when 936 => pixel <= "111111";
      when 937 => pixel <= "000000";
      when 938 => pixel <= "000000";
      when 939 => pixel <= "111111";
      when 940 => pixel <= "111111";
      when 941 => pixel <= "111111";
      when 942 => pixel <= "111111";
      when 943 => pixel <= "111111";
      when 944 => pixel <= "111111";
      when 945 => pixel <= "111111";
      when 946 => pixel <= "111111";
      when 947 => pixel <= "111111";
      when 948 => pixel <= "000000";
      when 949 => pixel <= "000000";
      when 950 => pixel <= "111111";
      when 951 => pixel <= "111111";
      when 952 => pixel <= "111111";
      when 953 => pixel <= "000000";
      when 954 => pixel <= "000000";
      when 955 => pixel <= "111111";
      when 956 => pixel <= "111111";
      when 957 => pixel <= "111111";
      when 958 => pixel <= "111111";
      when 959 => pixel <= "111111";
      when 960 => pixel <= "111111";
      when 961 => pixel <= "111111";
      when 962 => pixel <= "111111";
      when 963 => pixel <= "111111";
      when 964 => pixel <= "000000";
      when 965 => pixel <= "000000";
      when 966 => pixel <= "111111";
      when 967 => pixel <= "111111";
      when 968 => pixel <= "111111";
      when 969 => pixel <= "000000";
      when 970 => pixel <= "000000";
      when 971 => pixel <= "111111";
      when 972 => pixel <= "111111";
      when 973 => pixel <= "111111";
      when 974 => pixel <= "111111";
      when 975 => pixel <= "111111";
      when 976 => pixel <= "111111";
      when 977 => pixel <= "111111";
      when 978 => pixel <= "111111";
      when 979 => pixel <= "111111";
      when 980 => pixel <= "111111";
      when 981 => pixel <= "111111";
      when 982 => pixel <= "111111";
      when 983 => pixel <= "000000";
      when 984 => pixel <= "000000";
      when 985 => pixel <= "111111";
      when 986 => pixel <= "111111";
      when 987 => pixel <= "111111";
      when 988 => pixel <= "111111";
      when 989 => pixel <= "111111";
      when 990 => pixel <= "111111";
      when 991 => pixel <= "111111";
      when 992 => pixel <= "111111";
      when 993 => pixel <= "111111";
      when 994 => pixel <= "111111";
      when 995 => pixel <= "111111";
      when 996 => pixel <= "111111";
      when 997 => pixel <= "111111";
      when 998 => pixel <= "111111";
      when 999 => pixel <= "111111";
      when 1000 => pixel <= "000000";
      when 1001 => pixel <= "000000";
      when 1002 => pixel <= "111111";
      when 1003 => pixel <= "111111";
      when 1004 => pixel <= "111111";
      when 1005 => pixel <= "111111";
      when 1006 => pixel <= "111111";
      when 1007 => pixel <= "111111";
      when 1008 => pixel <= "111111";
      when 1009 => pixel <= "111111";
      when 1010 => pixel <= "111111";
      when 1011 => pixel <= "111111";
      when 1012 => pixel <= "111111";
      when 1013 => pixel <= "111111";
      when 1014 => pixel <= "111111";
      when 1015 => pixel <= "111111";
      when 1016 => pixel <= "111111";
      when 1017 => pixel <= "000000";
      when 1018 => pixel <= "000000";
      when 1019 => pixel <= "111111";
      when 1020 => pixel <= "111111";
      when 1021 => pixel <= "111111";
      when 1022 => pixel <= "111111";
      when 1023 => pixel <= "111111";
      when 1024 => pixel <= "111111";
      when 1025 => pixel <= "111111";
      when 1026 => pixel <= "111111";
      when 1027 => pixel <= "111111";
      when 1028 => pixel <= "111111";
      when 1029 => pixel <= "000000";
      when 1030 => pixel <= "000000";
      when 1031 => pixel <= "111111";
      when 1032 => pixel <= "000000";
      when 1033 => pixel <= "000000";
      when 1034 => pixel <= "111111";
      when 1035 => pixel <= "111111";
      when 1036 => pixel <= "111111";
      when 1037 => pixel <= "111111";
      when 1038 => pixel <= "111111";
      when 1039 => pixel <= "111111";
      when 1040 => pixel <= "111111";
      when 1041 => pixel <= "111111";
      when 1042 => pixel <= "111111";
      when 1043 => pixel <= "111111";
      when 1044 => pixel <= "000000";
      when 1045 => pixel <= "000000";
      when 1046 => pixel <= "111111";
      when 1047 => pixel <= "111111";
      when 1048 => pixel <= "111111";
      when 1049 => pixel <= "111111";
      when 1050 => pixel <= "111111";
      when 1051 => pixel <= "111111";
      when 1052 => pixel <= "111111";
      when 1053 => pixel <= "111111";
      when 1054 => pixel <= "111111";
      when 1055 => pixel <= "111111";
      when 1056 => pixel <= "111111";
      when 1057 => pixel <= "111111";
      when 1058 => pixel <= "111111";
      when 1059 => pixel <= "111111";
      when 1060 => pixel <= "000000";
      when 1061 => pixel <= "000000";
      when 1062 => pixel <= "111111";
      when 1063 => pixel <= "111111";
      when 1064 => pixel <= "111111";
      when 1065 => pixel <= "111111";
      when 1066 => pixel <= "111111";
      when 1067 => pixel <= "111111";
      when 1068 => pixel <= "111111";
      when 1069 => pixel <= "111111";
      when 1070 => pixel <= "111111";
      when 1071 => pixel <= "111111";
      when 1072 => pixel <= "111111";
      when 1073 => pixel <= "111111";
      when 1074 => pixel <= "111111";
      when 1075 => pixel <= "111111";
      when 1076 => pixel <= "111111";
      when 1077 => pixel <= "111111";
      when 1078 => pixel <= "111111";
      when 1079 => pixel <= "111111";
      when 1080 => pixel <= "111111";
      when 1081 => pixel <= "000000";
      when 1082 => pixel <= "000000";
      when 1083 => pixel <= "111111";
      when 1084 => pixel <= "111111";
      when 1085 => pixel <= "111111";
      when 1086 => pixel <= "111111";
      when 1087 => pixel <= "111111";
      when 1088 => pixel <= "111111";
      when 1089 => pixel <= "111111";
      when 1090 => pixel <= "111111";
      when 1091 => pixel <= "111111";
      when 1092 => pixel <= "000000";
      when 1093 => pixel <= "000000";
      when 1094 => pixel <= "111111";
      when 1095 => pixel <= "111111";
      when 1096 => pixel <= "111111";
      when 1097 => pixel <= "000000";
      when 1098 => pixel <= "000000";
      when 1099 => pixel <= "111111";
      when 1100 => pixel <= "111111";
      when 1101 => pixel <= "111111";
      when 1102 => pixel <= "111111";
      when 1103 => pixel <= "111111";
      when 1104 => pixel <= "111111";
      when 1105 => pixel <= "111111";
      when 1106 => pixel <= "111111";
      when 1107 => pixel <= "111111";
      when 1108 => pixel <= "000000";
      when 1109 => pixel <= "000000";
      when 1110 => pixel <= "111111";
      when 1111 => pixel <= "111111";
      when 1112 => pixel <= "111111";
      when 1113 => pixel <= "000000";
      when 1114 => pixel <= "000000";
      when 1115 => pixel <= "111111";
      when 1116 => pixel <= "111111";
      when 1117 => pixel <= "111111";
      when 1118 => pixel <= "111111";
      when 1119 => pixel <= "111111";
      when 1120 => pixel <= "111111";
      when 1121 => pixel <= "111111";
      when 1122 => pixel <= "111111";
      when 1123 => pixel <= "111111";
      when 1124 => pixel <= "000000";
      when 1125 => pixel <= "000000";
      when 1126 => pixel <= "111111";
      when 1127 => pixel <= "000000";
      when 1128 => pixel <= "111111";
      when 1129 => pixel <= "000000";
      when 1130 => pixel <= "000000";
      when 1131 => pixel <= "111111";
      when 1132 => pixel <= "111111";
      when 1133 => pixel <= "111111";
      when 1134 => pixel <= "111111";
      when 1135 => pixel <= "111111";
      when 1136 => pixel <= "111111";
      when 1137 => pixel <= "111111";
      when 1138 => pixel <= "111111";
      when 1139 => pixel <= "111111";
      when 1140 => pixel <= "111111";
      when 1141 => pixel <= "111111";
      when 1142 => pixel <= "111111";
      when 1143 => pixel <= "000000";
      when 1144 => pixel <= "000000";
      when 1145 => pixel <= "111111";
      when 1146 => pixel <= "111111";
      when 1147 => pixel <= "111111";
      when 1148 => pixel <= "111111";
      when 1149 => pixel <= "111111";
      when 1150 => pixel <= "111111";
      when 1151 => pixel <= "111111";
      when 1152 => pixel <= "111111";
      when 1153 => pixel <= "111111";
      when 1154 => pixel <= "111111";
      when 1155 => pixel <= "111111";
      when 1156 => pixel <= "111111";
      when 1157 => pixel <= "111111";
      when 1158 => pixel <= "111111";
      when 1159 => pixel <= "000000";
      when 1160 => pixel <= "000000";
      when 1161 => pixel <= "111111";
      when 1162 => pixel <= "111111";
      when 1163 => pixel <= "111111";
      when 1164 => pixel <= "111111";
      when 1165 => pixel <= "111111";
      when 1166 => pixel <= "111111";
      when 1167 => pixel <= "111111";
      when 1168 => pixel <= "111111";
      when 1169 => pixel <= "111111";
      when 1170 => pixel <= "111111";
      when 1171 => pixel <= "111111";
      when 1172 => pixel <= "111111";
      when 1173 => pixel <= "111111";
      when 1174 => pixel <= "000000";
      when 1175 => pixel <= "000000";
      when 1176 => pixel <= "000000";
      when 1177 => pixel <= "000000";
      when 1178 => pixel <= "111111";
      when 1179 => pixel <= "111111";
      when 1180 => pixel <= "111111";
      when 1181 => pixel <= "111111";
      when 1182 => pixel <= "111111";
      when 1183 => pixel <= "111111";
      when 1184 => pixel <= "111111";
      when 1185 => pixel <= "111111";
      when 1186 => pixel <= "111111";
      when 1187 => pixel <= "111111";
      when 1188 => pixel <= "000000";
      when 1189 => pixel <= "000000";
      when 1190 => pixel <= "111111";
      when 1191 => pixel <= "111111";
      when 1192 => pixel <= "000000";
      when 1193 => pixel <= "000000";
      when 1194 => pixel <= "111111";
      when 1195 => pixel <= "111111";
      when 1196 => pixel <= "111111";
      when 1197 => pixel <= "111111";
      when 1198 => pixel <= "111111";
      when 1199 => pixel <= "111111";
      when 1200 => pixel <= "111111";
      when 1201 => pixel <= "111111";
      when 1202 => pixel <= "111111";
      when 1203 => pixel <= "111111";
      when 1204 => pixel <= "000000";
      when 1205 => pixel <= "000000";
      when 1206 => pixel <= "000000";
      when 1207 => pixel <= "000000";
      when 1208 => pixel <= "000000";
      when 1209 => pixel <= "000000";
      when 1210 => pixel <= "111111";
      when 1211 => pixel <= "111111";
      when 1212 => pixel <= "111111";
      when 1213 => pixel <= "111111";
      when 1214 => pixel <= "111111";
      when 1215 => pixel <= "111111";
      when 1216 => pixel <= "111111";
      when 1217 => pixel <= "111111";
      when 1218 => pixel <= "111111";
      when 1219 => pixel <= "111111";
      when 1220 => pixel <= "000000";
      when 1221 => pixel <= "000000";
      when 1222 => pixel <= "000000";
      when 1223 => pixel <= "000000";
      when 1224 => pixel <= "000000";
      when 1225 => pixel <= "000000";
      when 1226 => pixel <= "111111";
      when 1227 => pixel <= "111111";
      when 1228 => pixel <= "111111";
      when 1229 => pixel <= "111111";
      when 1230 => pixel <= "111111";
      when 1231 => pixel <= "111111";
      when 1232 => pixel <= "111111";
      when 1233 => pixel <= "111111";
      when 1234 => pixel <= "111111";
      when 1235 => pixel <= "111111";
      when 1236 => pixel <= "111111";
      when 1237 => pixel <= "111111";
      when 1238 => pixel <= "111111";
      when 1239 => pixel <= "111111";
      when 1240 => pixel <= "000000";
      when 1241 => pixel <= "000000";
      when 1242 => pixel <= "111111";
      when 1243 => pixel <= "111111";
      when 1244 => pixel <= "111111";
      when 1245 => pixel <= "111111";
      when 1246 => pixel <= "111111";
      when 1247 => pixel <= "111111";
      when 1248 => pixel <= "111111";
      when 1249 => pixel <= "111111";
      when 1250 => pixel <= "111111";
      when 1251 => pixel <= "111111";
      when 1252 => pixel <= "111111";
      when 1253 => pixel <= "000000";
      when 1254 => pixel <= "000000";
      when 1255 => pixel <= "000000";
      when 1256 => pixel <= "000000";
      when 1257 => pixel <= "000000";
      when 1258 => pixel <= "111111";
      when 1259 => pixel <= "111111";
      when 1260 => pixel <= "111111";
      when 1261 => pixel <= "111111";
      when 1262 => pixel <= "111111";
      when 1263 => pixel <= "111111";
      when 1264 => pixel <= "111111";
      when 1265 => pixel <= "111111";
      when 1266 => pixel <= "111111";
      when 1267 => pixel <= "111111";
      when 1268 => pixel <= "111111";
      when 1269 => pixel <= "000000";
      when 1270 => pixel <= "000000";
      when 1271 => pixel <= "000000";
      when 1272 => pixel <= "000000";
      when 1273 => pixel <= "000000";
      when 1274 => pixel <= "000000";
      when 1275 => pixel <= "111111";
      when 1276 => pixel <= "111111";
      when 1277 => pixel <= "111111";
      when 1278 => pixel <= "111111";
      when 1279 => pixel <= "111111";
      when 1280 => pixel <= "111111";
      when 1281 => pixel <= "111111";
      when 1282 => pixel <= "111111";
      when 1283 => pixel <= "111111";
      when 1284 => pixel <= "000000";
      when 1285 => pixel <= "000000";
      when 1286 => pixel <= "111111";
      when 1287 => pixel <= "000000";
      when 1288 => pixel <= "111111";
      when 1289 => pixel <= "000000";
      when 1290 => pixel <= "000000";
      when 1291 => pixel <= "111111";
      when 1292 => pixel <= "111111";
      when 1293 => pixel <= "111111";
      when 1294 => pixel <= "111111";
      when 1295 => pixel <= "111111";
      when 1296 => pixel <= "111111";
      when 1297 => pixel <= "111111";
      when 1298 => pixel <= "111111";
      when 1299 => pixel <= "111111";
      when 1300 => pixel <= "111111";
      when 1301 => pixel <= "111111";
      when 1302 => pixel <= "111111";
      when 1303 => pixel <= "000000";
      when 1304 => pixel <= "000000";
      when 1305 => pixel <= "111111";
      when 1306 => pixel <= "111111";
      when 1307 => pixel <= "111111";
      when 1308 => pixel <= "111111";
      when 1309 => pixel <= "111111";
      when 1310 => pixel <= "111111";
      when 1311 => pixel <= "111111";
      when 1312 => pixel <= "111111";
      when 1313 => pixel <= "111111";
      when 1314 => pixel <= "111111";
      when 1315 => pixel <= "111111";
      when 1316 => pixel <= "111111";
      when 1317 => pixel <= "111111";
      when 1318 => pixel <= "000000";
      when 1319 => pixel <= "000000";
      when 1320 => pixel <= "111111";
      when 1321 => pixel <= "111111";
      when 1322 => pixel <= "111111";
      when 1323 => pixel <= "111111";
      when 1324 => pixel <= "111111";
      when 1325 => pixel <= "111111";
      when 1326 => pixel <= "111111";
      when 1327 => pixel <= "111111";
      when 1328 => pixel <= "111111";
      when 1329 => pixel <= "111111";
      when 1330 => pixel <= "111111";
      when 1331 => pixel <= "111111";
      when 1332 => pixel <= "111111";
      when 1333 => pixel <= "111111";
      when 1334 => pixel <= "111111";
      when 1335 => pixel <= "111111";
      when 1336 => pixel <= "111111";
      when 1337 => pixel <= "000000";
      when 1338 => pixel <= "000000";
      when 1339 => pixel <= "111111";
      when 1340 => pixel <= "111111";
      when 1341 => pixel <= "111111";
      when 1342 => pixel <= "111111";
      when 1343 => pixel <= "111111";
      when 1344 => pixel <= "111111";
      when 1345 => pixel <= "111111";
      when 1346 => pixel <= "111111";
      when 1347 => pixel <= "111111";
      when 1348 => pixel <= "000000";
      when 1349 => pixel <= "000000";
      when 1350 => pixel <= "000000";
      when 1351 => pixel <= "000000";
      when 1352 => pixel <= "000000";
      when 1353 => pixel <= "000000";
      when 1354 => pixel <= "000000";
      when 1355 => pixel <= "111111";
      when 1356 => pixel <= "111111";
      when 1357 => pixel <= "111111";
      when 1358 => pixel <= "111111";
      when 1359 => pixel <= "111111";
      when 1360 => pixel <= "111111";
      when 1361 => pixel <= "111111";
      when 1362 => pixel <= "111111";
      when 1363 => pixel <= "111111";
      when 1364 => pixel <= "111111";
      when 1365 => pixel <= "111111";
      when 1366 => pixel <= "111111";
      when 1367 => pixel <= "111111";
      when 1368 => pixel <= "111111";
      when 1369 => pixel <= "000000";
      when 1370 => pixel <= "000000";
      when 1371 => pixel <= "111111";
      when 1372 => pixel <= "111111";
      when 1373 => pixel <= "111111";
      when 1374 => pixel <= "111111";
      when 1375 => pixel <= "111111";
      when 1376 => pixel <= "111111";
      when 1377 => pixel <= "111111";
      when 1378 => pixel <= "111111";
      when 1379 => pixel <= "111111";
      when 1380 => pixel <= "000000";
      when 1381 => pixel <= "000000";
      when 1382 => pixel <= "111111";
      when 1383 => pixel <= "111111";
      when 1384 => pixel <= "111111";
      when 1385 => pixel <= "000000";
      when 1386 => pixel <= "000000";
      when 1387 => pixel <= "111111";
      when 1388 => pixel <= "111111";
      when 1389 => pixel <= "111111";
      when 1390 => pixel <= "111111";
      when 1391 => pixel <= "111111";
      when 1392 => pixel <= "111111";
      when 1393 => pixel <= "111111";
      when 1394 => pixel <= "111111";
      when 1395 => pixel <= "111111";
      when 1396 => pixel <= "111111";
      when 1397 => pixel <= "111111";
      when 1398 => pixel <= "111111";
      when 1399 => pixel <= "000000";
      when 1400 => pixel <= "000000";
      when 1401 => pixel <= "111111";
      when 1402 => pixel <= "111111";
      when 1403 => pixel <= "111111";
      when 1404 => pixel <= "111111";
      when 1405 => pixel <= "111111";
      when 1406 => pixel <= "111111";
      when 1407 => pixel <= "111111";
      when 1408 => pixel <= "111111";
      when 1409 => pixel <= "111111";
      when 1410 => pixel <= "111111";
      when 1411 => pixel <= "111111";
      when 1412 => pixel <= "000000";
      when 1413 => pixel <= "000000";
      when 1414 => pixel <= "111111";
      when 1415 => pixel <= "111111";
      when 1416 => pixel <= "111111";
      when 1417 => pixel <= "000000";
      when 1418 => pixel <= "000000";
      when 1419 => pixel <= "111111";
      when 1420 => pixel <= "111111";
      when 1421 => pixel <= "111111";
      when 1422 => pixel <= "111111";
      when 1423 => pixel <= "111111";
      when 1424 => pixel <= "111111";
      when 1425 => pixel <= "111111";
      when 1426 => pixel <= "111111";
      when 1427 => pixel <= "111111";
      when 1428 => pixel <= "111111";
      when 1429 => pixel <= "111111";
      when 1430 => pixel <= "111111";
      when 1431 => pixel <= "111111";
      when 1432 => pixel <= "111111";
      when 1433 => pixel <= "000000";
      when 1434 => pixel <= "000000";
      when 1435 => pixel <= "111111";
      when 1436 => pixel <= "111111";
      when 1437 => pixel <= "111111";
      when 1438 => pixel <= "111111";
      when 1439 => pixel <= "111111";
      when 1440 => pixel <= "111111";
      when 1441 => pixel <= "111111";
      when 1442 => pixel <= "111111";
      when 1443 => pixel <= "111111";
      when 1444 => pixel <= "000000";
      when 1445 => pixel <= "000000";
      when 1446 => pixel <= "111111";
      when 1447 => pixel <= "111111";
      when 1448 => pixel <= "111111";
      when 1449 => pixel <= "000000";
      when 1450 => pixel <= "000000";
      when 1451 => pixel <= "111111";
      when 1452 => pixel <= "111111";
      when 1453 => pixel <= "111111";
      when 1454 => pixel <= "111111";
      when 1455 => pixel <= "111111";
      when 1456 => pixel <= "111111";
      when 1457 => pixel <= "111111";
      when 1458 => pixel <= "111111";
      when 1459 => pixel <= "111111";
      when 1460 => pixel <= "111111";
      when 1461 => pixel <= "111111";
      when 1462 => pixel <= "111111";
      when 1463 => pixel <= "000000";
      when 1464 => pixel <= "000000";
      when 1465 => pixel <= "111111";
      when 1466 => pixel <= "111111";
      when 1467 => pixel <= "111111";
      when 1468 => pixel <= "111111";
      when 1469 => pixel <= "111111";
      when 1470 => pixel <= "111111";
      when 1471 => pixel <= "111111";
      when 1472 => pixel <= "111111";
      when 1473 => pixel <= "111111";
      when 1474 => pixel <= "111111";
      when 1475 => pixel <= "111111";
      when 1476 => pixel <= "111111";
      when 1477 => pixel <= "000000";
      when 1478 => pixel <= "000000";
      when 1479 => pixel <= "111111";
      when 1480 => pixel <= "111111";
      when 1481 => pixel <= "111111";
      when 1482 => pixel <= "111111";
      when 1483 => pixel <= "111111";
      when 1484 => pixel <= "111111";
      when 1485 => pixel <= "111111";
      when 1486 => pixel <= "111111";
      when 1487 => pixel <= "111111";
      when 1488 => pixel <= "111111";
      when 1489 => pixel <= "111111";
      when 1490 => pixel <= "111111";
      when 1491 => pixel <= "111111";
      when 1492 => pixel <= "111111";
      when 1493 => pixel <= "111111";
      when 1494 => pixel <= "111111";
      when 1495 => pixel <= "111111";
      when 1496 => pixel <= "111111";
      when 1497 => pixel <= "000000";
      when 1498 => pixel <= "000000";
      when 1499 => pixel <= "111111";
      when 1500 => pixel <= "111111";
      when 1501 => pixel <= "111111";
      when 1502 => pixel <= "111111";
      when 1503 => pixel <= "111111";
      when 1504 => pixel <= "111111";
      when 1505 => pixel <= "111111";
      when 1506 => pixel <= "111111";
      when 1507 => pixel <= "111111";
      when 1508 => pixel <= "111111";
      when 1509 => pixel <= "111111";
      when 1510 => pixel <= "111111";
      when 1511 => pixel <= "111111";
      when 1512 => pixel <= "000000";
      when 1513 => pixel <= "000000";
      when 1514 => pixel <= "111111";
      when 1515 => pixel <= "111111";
      when 1516 => pixel <= "111111";
      when 1517 => pixel <= "111111";
      when 1518 => pixel <= "111111";
      when 1519 => pixel <= "111111";
      when 1520 => pixel <= "111111";
      when 1521 => pixel <= "111111";
      when 1522 => pixel <= "111111";
      when 1523 => pixel <= "111111";
      when 1524 => pixel <= "111111";
      when 1525 => pixel <= "111111";
      when 1526 => pixel <= "111111";
      when 1527 => pixel <= "111111";
      when 1528 => pixel <= "111111";
      when 1529 => pixel <= "000000";
      when 1530 => pixel <= "000000";
      when 1531 => pixel <= "111111";
      when 1532 => pixel <= "111111";
      when 1533 => pixel <= "111111";
      when 1534 => pixel <= "111111";
      when 1535 => pixel <= "111111";
      when 1536 => pixel <= "111111";
      when 1537 => pixel <= "111111";
      when 1538 => pixel <= "111111";
      when 1539 => pixel <= "111111";
      when 1540 => pixel <= "000000";
      when 1541 => pixel <= "000000";
      when 1542 => pixel <= "111111";
      when 1543 => pixel <= "111111";
      when 1544 => pixel <= "111111";
      when 1545 => pixel <= "000000";
      when 1546 => pixel <= "000000";
      when 1547 => pixel <= "111111";
      when 1548 => pixel <= "111111";
      when 1549 => pixel <= "111111";
      when 1550 => pixel <= "111111";
      when 1551 => pixel <= "111111";
      when 1552 => pixel <= "111111";
      when 1553 => pixel <= "111111";
      when 1554 => pixel <= "111111";
      when 1555 => pixel <= "111111";
      when 1556 => pixel <= "111111";
      when 1557 => pixel <= "111111";
      when 1558 => pixel <= "000000";
      when 1559 => pixel <= "000000";
      when 1560 => pixel <= "111111";
      when 1561 => pixel <= "111111";
      when 1562 => pixel <= "111111";
      when 1563 => pixel <= "111111";
      when 1564 => pixel <= "111111";
      when 1565 => pixel <= "111111";
      when 1566 => pixel <= "111111";
      when 1567 => pixel <= "111111";
      when 1568 => pixel <= "111111";
      when 1569 => pixel <= "111111";
      when 1570 => pixel <= "111111";
      when 1571 => pixel <= "111111";
      when 1572 => pixel <= "000000";
      when 1573 => pixel <= "000000";
      when 1574 => pixel <= "111111";
      when 1575 => pixel <= "111111";
      when 1576 => pixel <= "111111";
      when 1577 => pixel <= "000000";
      when 1578 => pixel <= "000000";
      when 1579 => pixel <= "111111";
      when 1580 => pixel <= "111111";
      when 1581 => pixel <= "111111";
      when 1582 => pixel <= "111111";
      when 1583 => pixel <= "111111";
      when 1584 => pixel <= "111111";
      when 1585 => pixel <= "111111";
      when 1586 => pixel <= "111111";
      when 1587 => pixel <= "111111";
      when 1588 => pixel <= "111111";
      when 1589 => pixel <= "111111";
      when 1590 => pixel <= "111111";
      when 1591 => pixel <= "111111";
      when 1592 => pixel <= "111111";
      when 1593 => pixel <= "000000";
      when 1594 => pixel <= "000000";
      when 1595 => pixel <= "111111";
      when 1596 => pixel <= "111111";
      when 1597 => pixel <= "111111";
      when 1598 => pixel <= "111111";
      when 1599 => pixel <= "111111";
      when 1600 => pixel <= "111111";
      when 1601 => pixel <= "111111";
      when 1602 => pixel <= "111111";
      when 1603 => pixel <= "111111";
      when 1604 => pixel <= "000000";
      when 1605 => pixel <= "000000";
      when 1606 => pixel <= "111111";
      when 1607 => pixel <= "111111";
      when 1608 => pixel <= "111111";
      when 1609 => pixel <= "000000";
      when 1610 => pixel <= "000000";
      when 1611 => pixel <= "111111";
      when 1612 => pixel <= "111111";
      when 1613 => pixel <= "111111";
      when 1614 => pixel <= "111111";
      when 1615 => pixel <= "111111";
      when 1616 => pixel <= "111111";
      when 1617 => pixel <= "111111";
      when 1618 => pixel <= "111111";
      when 1619 => pixel <= "111111";
      when 1620 => pixel <= "111111";
      when 1621 => pixel <= "111111";
      when 1622 => pixel <= "111111";
      when 1623 => pixel <= "000000";
      when 1624 => pixel <= "000000";
      when 1625 => pixel <= "111111";
      when 1626 => pixel <= "111111";
      when 1627 => pixel <= "111111";
      when 1628 => pixel <= "111111";
      when 1629 => pixel <= "111111";
      when 1630 => pixel <= "111111";
      when 1631 => pixel <= "111111";
      when 1632 => pixel <= "111111";
      when 1633 => pixel <= "111111";
      when 1634 => pixel <= "111111";
      when 1635 => pixel <= "111111";
      when 1636 => pixel <= "000000";
      when 1637 => pixel <= "000000";
      when 1638 => pixel <= "111111";
      when 1639 => pixel <= "111111";
      when 1640 => pixel <= "111111";
      when 1641 => pixel <= "111111";
      when 1642 => pixel <= "111111";
      when 1643 => pixel <= "111111";
      when 1644 => pixel <= "111111";
      when 1645 => pixel <= "111111";
      when 1646 => pixel <= "111111";
      when 1647 => pixel <= "111111";
      when 1648 => pixel <= "111111";
      when 1649 => pixel <= "111111";
      when 1650 => pixel <= "111111";
      when 1651 => pixel <= "111111";
      when 1652 => pixel <= "111111";
      when 1653 => pixel <= "111111";
      when 1654 => pixel <= "111111";
      when 1655 => pixel <= "111111";
      when 1656 => pixel <= "111111";
      when 1657 => pixel <= "000000";
      when 1658 => pixel <= "000000";
      when 1659 => pixel <= "111111";
      when 1660 => pixel <= "111111";
      when 1661 => pixel <= "111111";
      when 1662 => pixel <= "111111";
      when 1663 => pixel <= "111111";
      when 1664 => pixel <= "111111";
      when 1665 => pixel <= "111111";
      when 1666 => pixel <= "111111";
      when 1667 => pixel <= "111111";
      when 1668 => pixel <= "111111";
      when 1669 => pixel <= "111111";
      when 1670 => pixel <= "111111";
      when 1671 => pixel <= "111111";
      when 1672 => pixel <= "000000";
      when 1673 => pixel <= "000000";
      when 1674 => pixel <= "111111";
      when 1675 => pixel <= "111111";
      when 1676 => pixel <= "111111";
      when 1677 => pixel <= "111111";
      when 1678 => pixel <= "111111";
      when 1679 => pixel <= "111111";
      when 1680 => pixel <= "111111";
      when 1681 => pixel <= "111111";
      when 1682 => pixel <= "111111";
      when 1683 => pixel <= "111111";
      when 1684 => pixel <= "111111";
      when 1685 => pixel <= "111111";
      when 1686 => pixel <= "111111";
      when 1687 => pixel <= "111111";
      when 1688 => pixel <= "111111";
      when 1689 => pixel <= "000000";
      when 1690 => pixel <= "000000";
      when 1691 => pixel <= "111111";
      when 1692 => pixel <= "111111";
      when 1693 => pixel <= "111111";
      when 1694 => pixel <= "111111";
      when 1695 => pixel <= "111111";
      when 1696 => pixel <= "111111";
      when 1697 => pixel <= "111111";
      when 1698 => pixel <= "111111";
      when 1699 => pixel <= "111111";
      when 1700 => pixel <= "000000";
      when 1701 => pixel <= "000000";
      when 1702 => pixel <= "111111";
      when 1703 => pixel <= "111111";
      when 1704 => pixel <= "111111";
      when 1705 => pixel <= "000000";
      when 1706 => pixel <= "000000";
      when 1707 => pixel <= "111111";
      when 1708 => pixel <= "111111";
      when 1709 => pixel <= "111111";
      when 1710 => pixel <= "111111";
      when 1711 => pixel <= "111111";
      when 1712 => pixel <= "111111";
      when 1713 => pixel <= "111111";
      when 1714 => pixel <= "111111";
      when 1715 => pixel <= "111111";
      when 1716 => pixel <= "111111";
      when 1717 => pixel <= "111111";
      when 1718 => pixel <= "000000";
      when 1719 => pixel <= "000000";
      when 1720 => pixel <= "111111";
      when 1721 => pixel <= "111111";
      when 1722 => pixel <= "111111";
      when 1723 => pixel <= "111111";
      when 1724 => pixel <= "111111";
      when 1725 => pixel <= "111111";
      when 1726 => pixel <= "111111";
      when 1727 => pixel <= "111111";
      when 1728 => pixel <= "111111";
      when 1729 => pixel <= "111111";
      when 1730 => pixel <= "111111";
      when 1731 => pixel <= "111111";
      when 1732 => pixel <= "000000";
      when 1733 => pixel <= "000000";
      when 1734 => pixel <= "111111";
      when 1735 => pixel <= "111111";
      when 1736 => pixel <= "111111";
      when 1737 => pixel <= "000000";
      when 1738 => pixel <= "000000";
      when 1739 => pixel <= "111111";
      when 1740 => pixel <= "111111";
      when 1741 => pixel <= "111111";
      when 1742 => pixel <= "111111";
      when 1743 => pixel <= "111111";
      when 1744 => pixel <= "111111";
      when 1745 => pixel <= "111111";
      when 1746 => pixel <= "111111";
      when 1747 => pixel <= "111111";
      when 1748 => pixel <= "111111";
      when 1749 => pixel <= "111111";
      when 1750 => pixel <= "111111";
      when 1751 => pixel <= "111111";
      when 1752 => pixel <= "111111";
      when 1753 => pixel <= "000000";
      when 1754 => pixel <= "000000";
      when 1755 => pixel <= "111111";
      when 1756 => pixel <= "111111";
      when 1757 => pixel <= "111111";
      when 1758 => pixel <= "111111";
      when 1759 => pixel <= "111111";
      when 1760 => pixel <= "111111";
      when 1761 => pixel <= "111111";
      when 1762 => pixel <= "111111";
      when 1763 => pixel <= "111111";
      when 1764 => pixel <= "111111";
      when 1765 => pixel <= "000000";
      when 1766 => pixel <= "000000";
      when 1767 => pixel <= "111111";
      when 1768 => pixel <= "000000";
      when 1769 => pixel <= "000000";
      when 1770 => pixel <= "111111";
      when 1771 => pixel <= "111111";
      when 1772 => pixel <= "111111";
      when 1773 => pixel <= "111111";
      when 1774 => pixel <= "111111";
      when 1775 => pixel <= "111111";
      when 1776 => pixel <= "111111";
      when 1777 => pixel <= "111111";
      when 1778 => pixel <= "111111";
      when 1779 => pixel <= "111111";
      when 1780 => pixel <= "111111";
      when 1781 => pixel <= "111111";
      when 1782 => pixel <= "111111";
      when 1783 => pixel <= "000000";
      when 1784 => pixel <= "000000";
      when 1785 => pixel <= "111111";
      when 1786 => pixel <= "111111";
      when 1787 => pixel <= "111111";
      when 1788 => pixel <= "111111";
      when 1789 => pixel <= "111111";
      when 1790 => pixel <= "111111";
      when 1791 => pixel <= "111111";
      when 1792 => pixel <= "111111";
      when 1793 => pixel <= "111111";
      when 1794 => pixel <= "111111";
      when 1795 => pixel <= "111111";
      when 1796 => pixel <= "000000";
      when 1797 => pixel <= "000000";
      when 1798 => pixel <= "111111";
      when 1799 => pixel <= "111111";
      when 1800 => pixel <= "111111";
      when 1801 => pixel <= "000000";
      when 1802 => pixel <= "000000";
      when 1803 => pixel <= "111111";
      when 1804 => pixel <= "111111";
      when 1805 => pixel <= "111111";
      when 1806 => pixel <= "111111";
      when 1807 => pixel <= "111111";
      when 1808 => pixel <= "111111";
      when 1809 => pixel <= "111111";
      when 1810 => pixel <= "111111";
      when 1811 => pixel <= "111111";
      when 1812 => pixel <= "000000";
      when 1813 => pixel <= "000000";
      when 1814 => pixel <= "111111";
      when 1815 => pixel <= "111111";
      when 1816 => pixel <= "111111";
      when 1817 => pixel <= "000000";
      when 1818 => pixel <= "000000";
      when 1819 => pixel <= "111111";
      when 1820 => pixel <= "111111";
      when 1821 => pixel <= "111111";
      when 1822 => pixel <= "111111";
      when 1823 => pixel <= "111111";
      when 1824 => pixel <= "111111";
      when 1825 => pixel <= "111111";
      when 1826 => pixel <= "111111";
      when 1827 => pixel <= "111111";
      when 1828 => pixel <= "111111";
      when 1829 => pixel <= "111111";
      when 1830 => pixel <= "111111";
      when 1831 => pixel <= "111111";
      when 1832 => pixel <= "000000";
      when 1833 => pixel <= "000000";
      when 1834 => pixel <= "111111";
      when 1835 => pixel <= "111111";
      when 1836 => pixel <= "111111";
      when 1837 => pixel <= "111111";
      when 1838 => pixel <= "111111";
      when 1839 => pixel <= "111111";
      when 1840 => pixel <= "111111";
      when 1841 => pixel <= "111111";
      when 1842 => pixel <= "111111";
      when 1843 => pixel <= "111111";
      when 1844 => pixel <= "000000";
      when 1845 => pixel <= "000000";
      when 1846 => pixel <= "111111";
      when 1847 => pixel <= "111111";
      when 1848 => pixel <= "111111";
      when 1849 => pixel <= "000000";
      when 1850 => pixel <= "000000";
      when 1851 => pixel <= "111111";
      when 1852 => pixel <= "111111";
      when 1853 => pixel <= "111111";
      when 1854 => pixel <= "111111";
      when 1855 => pixel <= "111111";
      when 1856 => pixel <= "111111";
      when 1857 => pixel <= "111111";
      when 1858 => pixel <= "111111";
      when 1859 => pixel <= "111111";
      when 1860 => pixel <= "000000";
      when 1861 => pixel <= "000000";
      when 1862 => pixel <= "111111";
      when 1863 => pixel <= "111111";
      when 1864 => pixel <= "111111";
      when 1865 => pixel <= "000000";
      when 1866 => pixel <= "000000";
      when 1867 => pixel <= "111111";
      when 1868 => pixel <= "111111";
      when 1869 => pixel <= "111111";
      when 1870 => pixel <= "111111";
      when 1871 => pixel <= "111111";
      when 1872 => pixel <= "111111";
      when 1873 => pixel <= "111111";
      when 1874 => pixel <= "111111";
      when 1875 => pixel <= "111111";
      when 1876 => pixel <= "111111";
      when 1877 => pixel <= "111111";
      when 1878 => pixel <= "000000";
      when 1879 => pixel <= "000000";
      when 1880 => pixel <= "111111";
      when 1881 => pixel <= "111111";
      when 1882 => pixel <= "111111";
      when 1883 => pixel <= "111111";
      when 1884 => pixel <= "111111";
      when 1885 => pixel <= "111111";
      when 1886 => pixel <= "111111";
      when 1887 => pixel <= "111111";
      when 1888 => pixel <= "111111";
      when 1889 => pixel <= "111111";
      when 1890 => pixel <= "111111";
      when 1891 => pixel <= "111111";
      when 1892 => pixel <= "000000";
      when 1893 => pixel <= "000000";
      when 1894 => pixel <= "111111";
      when 1895 => pixel <= "111111";
      when 1896 => pixel <= "111111";
      when 1897 => pixel <= "000000";
      when 1898 => pixel <= "000000";
      when 1899 => pixel <= "111111";
      when 1900 => pixel <= "111111";
      when 1901 => pixel <= "111111";
      when 1902 => pixel <= "111111";
      when 1903 => pixel <= "111111";
      when 1904 => pixel <= "111111";
      when 1905 => pixel <= "111111";
      when 1906 => pixel <= "111111";
      when 1907 => pixel <= "111111";
      when 1908 => pixel <= "111111";
      when 1909 => pixel <= "111111";
      when 1910 => pixel <= "111111";
      when 1911 => pixel <= "111111";
      when 1912 => pixel <= "000000";
      when 1913 => pixel <= "000000";
      when 1914 => pixel <= "111111";
      when 1915 => pixel <= "111111";
      when 1916 => pixel <= "111111";
      when 1917 => pixel <= "111111";
      when 1918 => pixel <= "111111";
      when 1919 => pixel <= "111111";
      when 1920 => pixel <= "111111";
      when 1921 => pixel <= "111111";
      when 1922 => pixel <= "111111";
      when 1923 => pixel <= "111111";
      when 1924 => pixel <= "111111";
      when 1925 => pixel <= "111111";
      when 1926 => pixel <= "000000";
      when 1927 => pixel <= "000000";
      when 1928 => pixel <= "000000";
      when 1929 => pixel <= "111111";
      when 1930 => pixel <= "111111";
      when 1931 => pixel <= "111111";
      when 1932 => pixel <= "111111";
      when 1933 => pixel <= "111111";
      when 1934 => pixel <= "111111";
      when 1935 => pixel <= "111111";
      when 1936 => pixel <= "111111";
      when 1937 => pixel <= "111111";
      when 1938 => pixel <= "111111";
      when 1939 => pixel <= "111111";
      when 1940 => pixel <= "111111";
      when 1941 => pixel <= "000000";
      when 1942 => pixel <= "000000";
      when 1943 => pixel <= "000000";
      when 1944 => pixel <= "000000";
      when 1945 => pixel <= "000000";
      when 1946 => pixel <= "000000";
      when 1947 => pixel <= "111111";
      when 1948 => pixel <= "111111";
      when 1949 => pixel <= "111111";
      when 1950 => pixel <= "111111";
      when 1951 => pixel <= "111111";
      when 1952 => pixel <= "111111";
      when 1953 => pixel <= "111111";
      when 1954 => pixel <= "111111";
      when 1955 => pixel <= "111111";
      when 1956 => pixel <= "000000";
      when 1957 => pixel <= "000000";
      when 1958 => pixel <= "000000";
      when 1959 => pixel <= "000000";
      when 1960 => pixel <= "000000";
      when 1961 => pixel <= "000000";
      when 1962 => pixel <= "000000";
      when 1963 => pixel <= "111111";
      when 1964 => pixel <= "111111";
      when 1965 => pixel <= "111111";
      when 1966 => pixel <= "111111";
      when 1967 => pixel <= "111111";
      when 1968 => pixel <= "111111";
      when 1969 => pixel <= "111111";
      when 1970 => pixel <= "111111";
      when 1971 => pixel <= "111111";
      when 1972 => pixel <= "111111";
      when 1973 => pixel <= "000000";
      when 1974 => pixel <= "000000";
      when 1975 => pixel <= "000000";
      when 1976 => pixel <= "000000";
      when 1977 => pixel <= "000000";
      when 1978 => pixel <= "111111";
      when 1979 => pixel <= "111111";
      when 1980 => pixel <= "111111";
      when 1981 => pixel <= "111111";
      when 1982 => pixel <= "111111";
      when 1983 => pixel <= "111111";
      when 1984 => pixel <= "111111";
      when 1985 => pixel <= "111111";
      when 1986 => pixel <= "111111";
      when 1987 => pixel <= "111111";
      when 1988 => pixel <= "111111";
      when 1989 => pixel <= "111111";
      when 1990 => pixel <= "111111";
      when 1991 => pixel <= "000000";
      when 1992 => pixel <= "000000";
      when 1993 => pixel <= "000000";
      when 1994 => pixel <= "000000";
      when 1995 => pixel <= "111111";
      when 1996 => pixel <= "111111";
      when 1997 => pixel <= "111111";
      when 1998 => pixel <= "111111";
      when 1999 => pixel <= "111111";
      when 2000 => pixel <= "111111";
      when 2001 => pixel <= "111111";
      when 2002 => pixel <= "111111";
      when 2003 => pixel <= "111111";
      when 2004 => pixel <= "111111";
      when 2005 => pixel <= "000000";
      when 2006 => pixel <= "000000";
      when 2007 => pixel <= "000000";
      when 2008 => pixel <= "000000";
      when 2009 => pixel <= "000000";
      when 2010 => pixel <= "111111";
      when 2011 => pixel <= "111111";
      when 2012 => pixel <= "111111";
      when 2013 => pixel <= "111111";
      when 2014 => pixel <= "111111";
      when 2015 => pixel <= "111111";
      when 2016 => pixel <= "111111";
      when 2017 => pixel <= "111111";
      when 2018 => pixel <= "111111";
      when 2019 => pixel <= "111111";
      when 2020 => pixel <= "111111";
      when 2021 => pixel <= "000000";
      when 2022 => pixel <= "000000";
      when 2023 => pixel <= "000000";
      when 2024 => pixel <= "000000";
      when 2025 => pixel <= "000000";
      when 2026 => pixel <= "111111";
      when 2027 => pixel <= "111111";
      when 2028 => pixel <= "111111";
      when 2029 => pixel <= "111111";
      when 2030 => pixel <= "111111";
      when 2031 => pixel <= "111111";
      when 2032 => pixel <= "111111";
      when 2033 => pixel <= "111111";
      when 2034 => pixel <= "111111";
      when 2035 => pixel <= "111111";
      when 2036 => pixel <= "111111";
      when 2037 => pixel <= "111111";
      when 2038 => pixel <= "000000";
      when 2039 => pixel <= "000000";
      when 2040 => pixel <= "111111";
      when 2041 => pixel <= "111111";
      when 2042 => pixel <= "111111";
      when 2043 => pixel <= "111111";
      when 2044 => pixel <= "111111";
      when 2045 => pixel <= "111111";
      when 2046 => pixel <= "111111";
      when 2047 => pixel <= "111111";
      when 2048 => pixel <= "111111";
      when 2049 => pixel <= "111111";
      when 2050 => pixel <= "111111";
      when 2051 => pixel <= "111111";
      when 2052 => pixel <= "111111";
      when 2053 => pixel <= "000000";
      when 2054 => pixel <= "000000";
      when 2055 => pixel <= "000000";
      when 2056 => pixel <= "000000";
      when 2057 => pixel <= "000000";
      when 2058 => pixel <= "111111";
      when 2059 => pixel <= "111111";
      when 2060 => pixel <= "111111";
      when 2061 => pixel <= "111111";
      when 2062 => pixel <= "111111";
      when 2063 => pixel <= "111111";
      when 2064 => pixel <= "111111";
      when 2065 => pixel <= "111111";
      when 2066 => pixel <= "111111";
      when 2067 => pixel <= "111111";
      when 2068 => pixel <= "111111";
      when 2069 => pixel <= "000000";
      when 2070 => pixel <= "000000";
      when 2071 => pixel <= "000000";
      when 2072 => pixel <= "000000";
      when 2073 => pixel <= "111111";
      when 2074 => pixel <= "111111";
      when 2075 => pixel <= "111111";
      when 2076 => pixel <= "111111";
      when 2077 => pixel <= "111111";
      when 2078 => pixel <= "111111";
      when 2079 => pixel <= "111111";
      when 2080 => pixel <= "111111";
      when 2081 => pixel <= "111111";
      when 2082 => pixel <= "111111";
      when 2083 => pixel <= "111111";
      when 2084 => pixel <= "111111";
      when 2085 => pixel <= "111111";
      when 2086 => pixel <= "111111";
      when 2087 => pixel <= "111111";
      when 2088 => pixel <= "111111";
      when 2089 => pixel <= "111111";
      when 2090 => pixel <= "111111";
      when 2091 => pixel <= "111111";
      when 2092 => pixel <= "111111";
      when 2093 => pixel <= "111111";
      when 2094 => pixel <= "111111";
      when 2095 => pixel <= "111111";
      when 2096 => pixel <= "111111";
      when 2097 => pixel <= "111111";
      when 2098 => pixel <= "111111";
      when 2099 => pixel <= "111111";
      when 2100 => pixel <= "111111";
      when 2101 => pixel <= "111111";
      when 2102 => pixel <= "111111";
      when 2103 => pixel <= "111111";
      when 2104 => pixel <= "111111";
      when 2105 => pixel <= "111111";
      when 2106 => pixel <= "111111";
      when 2107 => pixel <= "111111";
      when 2108 => pixel <= "111111";
      when 2109 => pixel <= "111111";
      when 2110 => pixel <= "111111";
      when 2111 => pixel <= "111111";
      when 2112 => pixel <= "111111";
      when 2113 => pixel <= "111111";
      when 2114 => pixel <= "111111";
      when 2115 => pixel <= "111111";
      when 2116 => pixel <= "111111";
      when 2117 => pixel <= "111111";
      when 2118 => pixel <= "111111";
      when 2119 => pixel <= "111111";
      when 2120 => pixel <= "111111";
      when 2121 => pixel <= "111111";
      when 2122 => pixel <= "111111";
      when 2123 => pixel <= "111111";
      when 2124 => pixel <= "111111";
      when 2125 => pixel <= "111111";
      when 2126 => pixel <= "111111";
      when 2127 => pixel <= "111111";
      when 2128 => pixel <= "111111";
      when 2129 => pixel <= "111111";
      when 2130 => pixel <= "111111";
      when 2131 => pixel <= "111111";
      when 2132 => pixel <= "111111";
      when 2133 => pixel <= "111111";
      when 2134 => pixel <= "111111";
      when 2135 => pixel <= "111111";
      when 2136 => pixel <= "111111";
      when 2137 => pixel <= "111111";
      when 2138 => pixel <= "111111";
      when 2139 => pixel <= "111111";
      when 2140 => pixel <= "111111";
      when 2141 => pixel <= "111111";
      when 2142 => pixel <= "111111";
      when 2143 => pixel <= "111111";
      when 2144 => pixel <= "111111";
      when 2145 => pixel <= "111111";
      when 2146 => pixel <= "111111";
      when 2147 => pixel <= "111111";
      when 2148 => pixel <= "111111";
      when 2149 => pixel <= "111111";
      when 2150 => pixel <= "111111";
      when 2151 => pixel <= "111111";
      when 2152 => pixel <= "111111";
      when 2153 => pixel <= "111111";
      when 2154 => pixel <= "111111";
      when 2155 => pixel <= "111111";
      when 2156 => pixel <= "111111";
      when 2157 => pixel <= "111111";
      when 2158 => pixel <= "111111";
      when 2159 => pixel <= "111111";
      when 2160 => pixel <= "111111";
      when 2161 => pixel <= "111111";
      when 2162 => pixel <= "111111";
      when 2163 => pixel <= "111111";
      when 2164 => pixel <= "111111";
      when 2165 => pixel <= "111111";
      when 2166 => pixel <= "111111";
      when 2167 => pixel <= "111111";
      when 2168 => pixel <= "111111";
      when 2169 => pixel <= "111111";
      when 2170 => pixel <= "111111";
      when 2171 => pixel <= "111111";
      when 2172 => pixel <= "111111";
      when 2173 => pixel <= "111111";
      when 2174 => pixel <= "111111";
      when 2175 => pixel <= "111111";
      when 2176 => pixel <= "111111";
      when 2177 => pixel <= "111111";
      when 2178 => pixel <= "111111";
      when 2179 => pixel <= "111111";
      when 2180 => pixel <= "111111";
      when 2181 => pixel <= "111111";
      when 2182 => pixel <= "111111";
      when 2183 => pixel <= "111111";
      when 2184 => pixel <= "111111";
      when 2185 => pixel <= "111111";
      when 2186 => pixel <= "111111";
      when 2187 => pixel <= "111111";
      when 2188 => pixel <= "111111";
      when 2189 => pixel <= "111111";
      when 2190 => pixel <= "111111";
      when 2191 => pixel <= "111111";
      when 2192 => pixel <= "111111";
      when 2193 => pixel <= "111111";
      when 2194 => pixel <= "111111";
      when 2195 => pixel <= "111111";
      when 2196 => pixel <= "111111";
      when 2197 => pixel <= "111111";
      when 2198 => pixel <= "111111";
      when 2199 => pixel <= "111111";
      when 2200 => pixel <= "111111";
      when 2201 => pixel <= "111111";
      when 2202 => pixel <= "111111";
      when 2203 => pixel <= "111111";
      when 2204 => pixel <= "111111";
      when 2205 => pixel <= "111111";
      when 2206 => pixel <= "111111";
      when 2207 => pixel <= "111111";
      when 2208 => pixel <= "111111";
      when 2209 => pixel <= "111111";
      when 2210 => pixel <= "111111";
      when 2211 => pixel <= "111111";
      when 2212 => pixel <= "111111";
      when 2213 => pixel <= "111111";
      when 2214 => pixel <= "111111";
      when 2215 => pixel <= "111111";
      when 2216 => pixel <= "111111";
      when 2217 => pixel <= "111111";
      when 2218 => pixel <= "111111";
      when 2219 => pixel <= "111111";
      when 2220 => pixel <= "111111";
      when 2221 => pixel <= "111111";
      when 2222 => pixel <= "111111";
      when 2223 => pixel <= "111111";
      when 2224 => pixel <= "111111";
      when 2225 => pixel <= "111111";
      when 2226 => pixel <= "111111";
      when 2227 => pixel <= "111111";
      when 2228 => pixel <= "111111";
      when 2229 => pixel <= "111111";
      when 2230 => pixel <= "111111";
      when 2231 => pixel <= "111111";
      when 2232 => pixel <= "111111";
      when 2233 => pixel <= "111111";
      when 2234 => pixel <= "111111";
      when 2235 => pixel <= "111111";
      when 2236 => pixel <= "111111";
      when 2237 => pixel <= "111111";
      when 2238 => pixel <= "111111";
      when 2239 => pixel <= "111111";
      when 2240 => pixel <= "111111";
      when 2241 => pixel <= "111111";
      when 2242 => pixel <= "111111";
      when 2243 => pixel <= "111111";
      when 2244 => pixel <= "111111";
      when 2245 => pixel <= "111111";
      when 2246 => pixel <= "111111";
      when 2247 => pixel <= "111111";
      when 2248 => pixel <= "111111";
      when 2249 => pixel <= "111111";
      when 2250 => pixel <= "111111";
      when 2251 => pixel <= "111111";
      when 2252 => pixel <= "111111";
      when 2253 => pixel <= "111111";
      when 2254 => pixel <= "111111";
      when 2255 => pixel <= "111111";
      when 2256 => pixel <= "111111";
      when 2257 => pixel <= "111111";
      when 2258 => pixel <= "111111";
      when 2259 => pixel <= "111111";
      when 2260 => pixel <= "111111";
      when 2261 => pixel <= "111111";
      when 2262 => pixel <= "111111";
      when 2263 => pixel <= "111111";
      when 2264 => pixel <= "111111";
      when 2265 => pixel <= "111111";
      when 2266 => pixel <= "111111";
      when 2267 => pixel <= "111111";
      when 2268 => pixel <= "111111";
      when 2269 => pixel <= "111111";
      when 2270 => pixel <= "111111";
      when 2271 => pixel <= "111111";
      when 2272 => pixel <= "111111";
      when 2273 => pixel <= "111111";
      when 2274 => pixel <= "111111";
      when 2275 => pixel <= "111111";
      when 2276 => pixel <= "111111";
      when 2277 => pixel <= "111111";
      when 2278 => pixel <= "111111";
      when 2279 => pixel <= "111111";
      when 2280 => pixel <= "111111";
      when 2281 => pixel <= "111111";
      when 2282 => pixel <= "111111";
      when 2283 => pixel <= "111111";
      when 2284 => pixel <= "111111";
      when 2285 => pixel <= "111111";
      when 2286 => pixel <= "111111";
      when 2287 => pixel <= "111111";
      when 2288 => pixel <= "111111";
      when 2289 => pixel <= "111111";
      when 2290 => pixel <= "111111";
      when 2291 => pixel <= "111111";
      when 2292 => pixel <= "111111";
      when 2293 => pixel <= "111111";
      when 2294 => pixel <= "111111";
      when 2295 => pixel <= "111111";
      when 2296 => pixel <= "111111";
      when 2297 => pixel <= "111111";
      when 2298 => pixel <= "111111";
      when 2299 => pixel <= "111111";
      when 2300 => pixel <= "111111";
      when 2301 => pixel <= "111111";
      when 2302 => pixel <= "111111";
      when 2303 => pixel <= "111111";
      when 2304 => pixel <= "111111";
      when 2305 => pixel <= "111111";
      when 2306 => pixel <= "111111";
      when 2307 => pixel <= "111111";
      when 2308 => pixel <= "111111";
      when 2309 => pixel <= "111111";
      when 2310 => pixel <= "111111";
      when 2311 => pixel <= "111111";
      when 2312 => pixel <= "111111";
      when 2313 => pixel <= "111111";
      when 2314 => pixel <= "111111";
      when 2315 => pixel <= "111111";
      when 2316 => pixel <= "111111";
      when 2317 => pixel <= "111111";
      when 2318 => pixel <= "111111";
      when 2319 => pixel <= "111111";
      when 2320 => pixel <= "111111";
      when 2321 => pixel <= "111111";
      when 2322 => pixel <= "111111";
      when 2323 => pixel <= "111111";
      when 2324 => pixel <= "111111";
      when 2325 => pixel <= "111111";
      when 2326 => pixel <= "111111";
      when 2327 => pixel <= "111111";
      when 2328 => pixel <= "111111";
      when 2329 => pixel <= "111111";
      when 2330 => pixel <= "111111";
      when 2331 => pixel <= "111111";
      when 2332 => pixel <= "111111";
      when 2333 => pixel <= "111111";
      when 2334 => pixel <= "111111";
      when 2335 => pixel <= "111111";
      when 2336 => pixel <= "111111";
      when 2337 => pixel <= "111111";
      when 2338 => pixel <= "111111";
      when 2339 => pixel <= "111111";
      when 2340 => pixel <= "111111";
      when 2341 => pixel <= "111111";
      when 2342 => pixel <= "111111";
      when 2343 => pixel <= "111111";
      when 2344 => pixel <= "111111";
      when 2345 => pixel <= "111111";
      when 2346 => pixel <= "111111";
      when 2347 => pixel <= "111111";
      when 2348 => pixel <= "111111";
      when 2349 => pixel <= "111111";
      when 2350 => pixel <= "111111";
      when 2351 => pixel <= "111111";
      when 2352 => pixel <= "111111";
      when 2353 => pixel <= "111111";
      when 2354 => pixel <= "111111";
      when 2355 => pixel <= "111111";
      when 2356 => pixel <= "111111";
      when 2357 => pixel <= "111111";
      when 2358 => pixel <= "111111";
      when 2359 => pixel <= "111111";
      when 2360 => pixel <= "111111";
      when 2361 => pixel <= "111111";
      when 2362 => pixel <= "111111";
      when 2363 => pixel <= "111111";
      when 2364 => pixel <= "111111";
      when 2365 => pixel <= "111111";
      when 2366 => pixel <= "111111";
      when 2367 => pixel <= "111111";
      when 2368 => pixel <= "111111";
      when 2369 => pixel <= "111111";
      when 2370 => pixel <= "111111";
      when 2371 => pixel <= "111111";
      when 2372 => pixel <= "111111";
      when 2373 => pixel <= "111111";
      when 2374 => pixel <= "111111";
      when 2375 => pixel <= "111111";
      when 2376 => pixel <= "111111";
      when 2377 => pixel <= "111111";
      when 2378 => pixel <= "111111";
      when 2379 => pixel <= "111111";
      when 2380 => pixel <= "111111";
      when 2381 => pixel <= "111111";
      when 2382 => pixel <= "111111";
      when 2383 => pixel <= "111111";
      when 2384 => pixel <= "111111";
      when 2385 => pixel <= "111111";
      when 2386 => pixel <= "111111";
      when 2387 => pixel <= "111111";
      when 2388 => pixel <= "111111";
      when 2389 => pixel <= "111111";
      when 2390 => pixel <= "111111";
      when 2391 => pixel <= "111111";
      when 2392 => pixel <= "111111";
      when 2393 => pixel <= "111111";
      when 2394 => pixel <= "111111";
      when 2395 => pixel <= "111111";
      when 2396 => pixel <= "111111";
      when 2397 => pixel <= "111111";
      when 2398 => pixel <= "111111";
      when 2399 => pixel <= "111111";
      when 2400 => pixel <= "111111";
      when 2401 => pixel <= "111111";
      when 2402 => pixel <= "111111";
      when 2403 => pixel <= "111111";
      when 2404 => pixel <= "111111";
      when 2405 => pixel <= "111111";
      when 2406 => pixel <= "111111";
      when 2407 => pixel <= "111111";
      when 2408 => pixel <= "111111";
      when 2409 => pixel <= "111111";
      when 2410 => pixel <= "111111";
      when 2411 => pixel <= "111111";
      when 2412 => pixel <= "111111";
      when 2413 => pixel <= "111111";
      when 2414 => pixel <= "111111";
      when 2415 => pixel <= "111111";
      when 2416 => pixel <= "111111";
      when 2417 => pixel <= "111111";
      when 2418 => pixel <= "111111";
      when 2419 => pixel <= "111111";
      when 2420 => pixel <= "111111";
      when 2421 => pixel <= "111111";
      when 2422 => pixel <= "111111";
      when 2423 => pixel <= "111111";
      when 2424 => pixel <= "111111";
      when 2425 => pixel <= "111111";
      when 2426 => pixel <= "111111";
      when 2427 => pixel <= "111111";
      when 2428 => pixel <= "111111";
      when 2429 => pixel <= "111111";
      when 2430 => pixel <= "111111";
      when 2431 => pixel <= "111111";
      when 2432 => pixel <= "111111";
      when 2433 => pixel <= "111111";
      when 2434 => pixel <= "111111";
      when 2435 => pixel <= "111111";
      when 2436 => pixel <= "111111";
      when 2437 => pixel <= "111111";
      when 2438 => pixel <= "111111";
      when 2439 => pixel <= "111111";
      when 2440 => pixel <= "111111";
      when 2441 => pixel <= "111111";
      when 2442 => pixel <= "111111";
      when 2443 => pixel <= "111111";
      when 2444 => pixel <= "111111";
      when 2445 => pixel <= "111111";
      when 2446 => pixel <= "111111";
      when 2447 => pixel <= "111111";
      when 2448 => pixel <= "111111";
      when 2449 => pixel <= "111111";
      when 2450 => pixel <= "111111";
      when 2451 => pixel <= "111111";
      when 2452 => pixel <= "111111";
      when 2453 => pixel <= "111111";
      when 2454 => pixel <= "111111";
      when 2455 => pixel <= "111111";
      when 2456 => pixel <= "111111";
      when 2457 => pixel <= "111111";
      when 2458 => pixel <= "111111";
      when 2459 => pixel <= "111111";
      when 2460 => pixel <= "111111";
      when 2461 => pixel <= "111111";
      when 2462 => pixel <= "111111";
      when 2463 => pixel <= "111111";
      when 2464 => pixel <= "111111";
      when 2465 => pixel <= "111111";
      when 2466 => pixel <= "111111";
      when 2467 => pixel <= "111111";
      when 2468 => pixel <= "111111";
      when 2469 => pixel <= "111111";
      when 2470 => pixel <= "111111";
      when 2471 => pixel <= "111111";
      when 2472 => pixel <= "111111";
      when 2473 => pixel <= "111111";
      when 2474 => pixel <= "111111";
      when 2475 => pixel <= "111111";
      when 2476 => pixel <= "111111";
      when 2477 => pixel <= "111111";
      when 2478 => pixel <= "111111";
      when 2479 => pixel <= "111111";
      when 2480 => pixel <= "111111";
      when 2481 => pixel <= "111111";
      when 2482 => pixel <= "111111";
      when 2483 => pixel <= "111111";
      when 2484 => pixel <= "111111";
      when 2485 => pixel <= "111111";
      when 2486 => pixel <= "111111";
      when 2487 => pixel <= "111111";
      when 2488 => pixel <= "111111";
      when 2489 => pixel <= "111111";
      when 2490 => pixel <= "111111";
      when 2491 => pixel <= "111111";
      when 2492 => pixel <= "111111";
      when 2493 => pixel <= "111111";
      when 2494 => pixel <= "111111";
      when 2495 => pixel <= "111111";
      when 2496 => pixel <= "111111";
      when 2497 => pixel <= "111111";
      when 2498 => pixel <= "111111";
      when 2499 => pixel <= "111111";
      when 2500 => pixel <= "111111";
      when 2501 => pixel <= "111111";
      when 2502 => pixel <= "111111";
      when 2503 => pixel <= "111111";
      when 2504 => pixel <= "111111";
      when 2505 => pixel <= "111111";
      when 2506 => pixel <= "111111";
      when 2507 => pixel <= "111111";
      when 2508 => pixel <= "111111";
      when 2509 => pixel <= "111111";
      when 2510 => pixel <= "111111";
      when 2511 => pixel <= "111111";
      when 2512 => pixel <= "111111";
      when 2513 => pixel <= "111111";
      when 2514 => pixel <= "111111";
      when 2515 => pixel <= "111111";
      when 2516 => pixel <= "111111";
      when 2517 => pixel <= "111111";
      when 2518 => pixel <= "111111";
      when 2519 => pixel <= "111111";
      when 2520 => pixel <= "111111";
      when 2521 => pixel <= "111111";
      when 2522 => pixel <= "111111";
      when 2523 => pixel <= "111111";
      when 2524 => pixel <= "111111";
      when 2525 => pixel <= "111111";
      when 2526 => pixel <= "111111";
      when 2527 => pixel <= "111111";
      when 2528 => pixel <= "111111";
      when 2529 => pixel <= "111111";
      when 2530 => pixel <= "111111";
      when 2531 => pixel <= "111111";
      when 2532 => pixel <= "111111";
      when 2533 => pixel <= "111111";
      when 2534 => pixel <= "111111";
      when 2535 => pixel <= "111111";
      when 2536 => pixel <= "111111";
      when 2537 => pixel <= "111111";
      when 2538 => pixel <= "111111";
      when 2539 => pixel <= "111111";
      when 2540 => pixel <= "111111";
      when 2541 => pixel <= "111111";
      when 2542 => pixel <= "111111";
      when 2543 => pixel <= "111111";
      when 2544 => pixel <= "111111";
      when 2545 => pixel <= "111111";
      when 2546 => pixel <= "111111";
      when 2547 => pixel <= "111111";
      when 2548 => pixel <= "111111";
      when 2549 => pixel <= "111111";
      when 2550 => pixel <= "111111";
      when 2551 => pixel <= "111111";
      when 2552 => pixel <= "111111";
      when 2553 => pixel <= "111111";
      when 2554 => pixel <= "111111";
      when 2555 => pixel <= "111111";
      when 2556 => pixel <= "111111";
      when 2557 => pixel <= "111111";
      when 2558 => pixel <= "111111";
      when 2559 => pixel <= "111111";
      when others => pixel <= (others => '0');
    end case;
  end process;
end;
